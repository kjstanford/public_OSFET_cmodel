** gc array model

.TEMP 25.0
.OPTION
+ ARTIST=2
+ INGOLD=2
+ PARHIER=LOCAL
+ PSF=2
+ ACCURATE=1
+ POST=2

.HDL "osfet_potential_based_compact_model_v0.va"
.INC "../model_card/rfet_params_v0.inc"
.INC "../model_card/wfet_params_v0.inc"

.PARAM vdd = 0.9
.PARAM vss = 0
.PARAM vpp = 1.2
.PARAM vnn = 0
.PARAM Rwwl = 100
.PARAM Cwwl = 1e-15
.PARAM Rwbl = 100
.PARAM Cwbl = 1e-15
.PARAM Rrwl = 100
.PARAM Crwl = 1e-15
.PARAM Rrbl = 100
.PARAM Crbl = 1e-15
.PARAM sim_time = 40e-9
.PARAM timestep = 1e-12
.SUBCKT wos_ros_gc wwl wbl rwl rbl sn

    xos wbl wwl sn osfet
    + W=W_write mu_eff=mu_eff_write Lch=Lch_write Cgch=Cgch_write Cpar=Cpar_write longVT=longVT_write alpha1=alpha1_write alpha2=alpha2_write meff=meff_write
    + rsd_mode=rsd_mode_write Rs0=Rs0_write Rd0=Rd0_write delta=delta_write rollVT=rollVT_write n0=n0_write nd=nd_write type=type_write

    xosr rbl sn rwl osfet
    + W=W_read mu_eff=mu_eff_read Lch=Lch_read Cgch=Cgch_read Cpar=Cpar_read longVT=longVT_read alpha1=alpha1_read alpha2=alpha2_read meff=meff_read
    + rsd_mode=rsd_mode_read Rs0=Rs0_read Rd0=Rd0_read delta=delta_read rollVT=rollVT_read n0=n0_read nd=nd_read type=type_read

.ENDS

.SUBCKT rc_unit rc_in rc_out R0=1e2 C0=1e-15

    r_unit rc_in rc_out R=R0
    c_unit rc_out 0 C=C0

.ENDS rc_unit
.DCVOLT sn_0_0 '0*vdd + 1*vss'
.DCVOLT sn_0_1 '0*vdd + 1*vss'
.DCVOLT sn_0_2 '0*vdd + 1*vss'
.DCVOLT sn_0_3 '0*vdd + 1*vss'
.DCVOLT sn_0_4 '0*vdd + 1*vss'
.DCVOLT sn_0_5 '0*vdd + 1*vss'
.DCVOLT sn_0_6 '0*vdd + 1*vss'
.DCVOLT sn_0_7 '0*vdd + 1*vss'
.DCVOLT sn_0_8 '0*vdd + 1*vss'
.DCVOLT sn_0_9 '0*vdd + 1*vss'
.DCVOLT sn_0_10 '0*vdd + 1*vss'
.DCVOLT sn_0_11 '0*vdd + 1*vss'
.DCVOLT sn_0_12 '0*vdd + 1*vss'
.DCVOLT sn_0_13 '0*vdd + 1*vss'
.DCVOLT sn_0_14 '0*vdd + 1*vss'
.DCVOLT sn_0_15 '0*vdd + 1*vss'
.DCVOLT sn_0_16 '0*vdd + 1*vss'
.DCVOLT sn_0_17 '0*vdd + 1*vss'
.DCVOLT sn_0_18 '0*vdd + 1*vss'
.DCVOLT sn_0_19 '0*vdd + 1*vss'
.DCVOLT sn_0_20 '0*vdd + 1*vss'
.DCVOLT sn_0_21 '0*vdd + 1*vss'
.DCVOLT sn_0_22 '0*vdd + 1*vss'
.DCVOLT sn_0_23 '0*vdd + 1*vss'
.DCVOLT sn_0_24 '0*vdd + 1*vss'
.DCVOLT sn_0_25 '0*vdd + 1*vss'
.DCVOLT sn_0_26 '0*vdd + 1*vss'
.DCVOLT sn_0_27 '0*vdd + 1*vss'
.DCVOLT sn_0_28 '0*vdd + 1*vss'
.DCVOLT sn_0_29 '0*vdd + 1*vss'
.DCVOLT sn_0_30 '0*vdd + 1*vss'
.DCVOLT sn_0_31 '0*vdd + 1*vss'
.DCVOLT sn_1_0 '0*vdd + 1*vss'
.DCVOLT sn_1_1 '0*vdd + 1*vss'
.DCVOLT sn_1_2 '0*vdd + 1*vss'
.DCVOLT sn_1_3 '0*vdd + 1*vss'
.DCVOLT sn_1_4 '0*vdd + 1*vss'
.DCVOLT sn_1_5 '0*vdd + 1*vss'
.DCVOLT sn_1_6 '0*vdd + 1*vss'
.DCVOLT sn_1_7 '0*vdd + 1*vss'
.DCVOLT sn_1_8 '0*vdd + 1*vss'
.DCVOLT sn_1_9 '0*vdd + 1*vss'
.DCVOLT sn_1_10 '0*vdd + 1*vss'
.DCVOLT sn_1_11 '0*vdd + 1*vss'
.DCVOLT sn_1_12 '0*vdd + 1*vss'
.DCVOLT sn_1_13 '0*vdd + 1*vss'
.DCVOLT sn_1_14 '0*vdd + 1*vss'
.DCVOLT sn_1_15 '0*vdd + 1*vss'
.DCVOLT sn_1_16 '0*vdd + 1*vss'
.DCVOLT sn_1_17 '0*vdd + 1*vss'
.DCVOLT sn_1_18 '0*vdd + 1*vss'
.DCVOLT sn_1_19 '0*vdd + 1*vss'
.DCVOLT sn_1_20 '0*vdd + 1*vss'
.DCVOLT sn_1_21 '0*vdd + 1*vss'
.DCVOLT sn_1_22 '0*vdd + 1*vss'
.DCVOLT sn_1_23 '0*vdd + 1*vss'
.DCVOLT sn_1_24 '0*vdd + 1*vss'
.DCVOLT sn_1_25 '0*vdd + 1*vss'
.DCVOLT sn_1_26 '0*vdd + 1*vss'
.DCVOLT sn_1_27 '0*vdd + 1*vss'
.DCVOLT sn_1_28 '0*vdd + 1*vss'
.DCVOLT sn_1_29 '0*vdd + 1*vss'
.DCVOLT sn_1_30 '0*vdd + 1*vss'
.DCVOLT sn_1_31 '0*vdd + 1*vss'
.DCVOLT sn_2_0 '0*vdd + 1*vss'
.DCVOLT sn_2_1 '0*vdd + 1*vss'
.DCVOLT sn_2_2 '0*vdd + 1*vss'
.DCVOLT sn_2_3 '0*vdd + 1*vss'
.DCVOLT sn_2_4 '0*vdd + 1*vss'
.DCVOLT sn_2_5 '0*vdd + 1*vss'
.DCVOLT sn_2_6 '0*vdd + 1*vss'
.DCVOLT sn_2_7 '0*vdd + 1*vss'
.DCVOLT sn_2_8 '0*vdd + 1*vss'
.DCVOLT sn_2_9 '0*vdd + 1*vss'
.DCVOLT sn_2_10 '0*vdd + 1*vss'
.DCVOLT sn_2_11 '0*vdd + 1*vss'
.DCVOLT sn_2_12 '0*vdd + 1*vss'
.DCVOLT sn_2_13 '0*vdd + 1*vss'
.DCVOLT sn_2_14 '0*vdd + 1*vss'
.DCVOLT sn_2_15 '0*vdd + 1*vss'
.DCVOLT sn_2_16 '0*vdd + 1*vss'
.DCVOLT sn_2_17 '0*vdd + 1*vss'
.DCVOLT sn_2_18 '0*vdd + 1*vss'
.DCVOLT sn_2_19 '0*vdd + 1*vss'
.DCVOLT sn_2_20 '0*vdd + 1*vss'
.DCVOLT sn_2_21 '0*vdd + 1*vss'
.DCVOLT sn_2_22 '0*vdd + 1*vss'
.DCVOLT sn_2_23 '0*vdd + 1*vss'
.DCVOLT sn_2_24 '0*vdd + 1*vss'
.DCVOLT sn_2_25 '0*vdd + 1*vss'
.DCVOLT sn_2_26 '0*vdd + 1*vss'
.DCVOLT sn_2_27 '0*vdd + 1*vss'
.DCVOLT sn_2_28 '0*vdd + 1*vss'
.DCVOLT sn_2_29 '0*vdd + 1*vss'
.DCVOLT sn_2_30 '0*vdd + 1*vss'
.DCVOLT sn_2_31 '0*vdd + 1*vss'
.DCVOLT sn_3_0 '0*vdd + 1*vss'
.DCVOLT sn_3_1 '0*vdd + 1*vss'
.DCVOLT sn_3_2 '0*vdd + 1*vss'
.DCVOLT sn_3_3 '0*vdd + 1*vss'
.DCVOLT sn_3_4 '0*vdd + 1*vss'
.DCVOLT sn_3_5 '0*vdd + 1*vss'
.DCVOLT sn_3_6 '0*vdd + 1*vss'
.DCVOLT sn_3_7 '0*vdd + 1*vss'
.DCVOLT sn_3_8 '0*vdd + 1*vss'
.DCVOLT sn_3_9 '0*vdd + 1*vss'
.DCVOLT sn_3_10 '0*vdd + 1*vss'
.DCVOLT sn_3_11 '0*vdd + 1*vss'
.DCVOLT sn_3_12 '0*vdd + 1*vss'
.DCVOLT sn_3_13 '0*vdd + 1*vss'
.DCVOLT sn_3_14 '0*vdd + 1*vss'
.DCVOLT sn_3_15 '0*vdd + 1*vss'
.DCVOLT sn_3_16 '0*vdd + 1*vss'
.DCVOLT sn_3_17 '0*vdd + 1*vss'
.DCVOLT sn_3_18 '0*vdd + 1*vss'
.DCVOLT sn_3_19 '0*vdd + 1*vss'
.DCVOLT sn_3_20 '0*vdd + 1*vss'
.DCVOLT sn_3_21 '0*vdd + 1*vss'
.DCVOLT sn_3_22 '0*vdd + 1*vss'
.DCVOLT sn_3_23 '0*vdd + 1*vss'
.DCVOLT sn_3_24 '0*vdd + 1*vss'
.DCVOLT sn_3_25 '0*vdd + 1*vss'
.DCVOLT sn_3_26 '0*vdd + 1*vss'
.DCVOLT sn_3_27 '0*vdd + 1*vss'
.DCVOLT sn_3_28 '0*vdd + 1*vss'
.DCVOLT sn_3_29 '0*vdd + 1*vss'
.DCVOLT sn_3_30 '0*vdd + 1*vss'
.DCVOLT sn_3_31 '0*vdd + 1*vss'
.DCVOLT sn_4_0 '0*vdd + 1*vss'
.DCVOLT sn_4_1 '0*vdd + 1*vss'
.DCVOLT sn_4_2 '0*vdd + 1*vss'
.DCVOLT sn_4_3 '0*vdd + 1*vss'
.DCVOLT sn_4_4 '0*vdd + 1*vss'
.DCVOLT sn_4_5 '0*vdd + 1*vss'
.DCVOLT sn_4_6 '0*vdd + 1*vss'
.DCVOLT sn_4_7 '0*vdd + 1*vss'
.DCVOLT sn_4_8 '0*vdd + 1*vss'
.DCVOLT sn_4_9 '0*vdd + 1*vss'
.DCVOLT sn_4_10 '0*vdd + 1*vss'
.DCVOLT sn_4_11 '0*vdd + 1*vss'
.DCVOLT sn_4_12 '0*vdd + 1*vss'
.DCVOLT sn_4_13 '0*vdd + 1*vss'
.DCVOLT sn_4_14 '0*vdd + 1*vss'
.DCVOLT sn_4_15 '0*vdd + 1*vss'
.DCVOLT sn_4_16 '0*vdd + 1*vss'
.DCVOLT sn_4_17 '0*vdd + 1*vss'
.DCVOLT sn_4_18 '0*vdd + 1*vss'
.DCVOLT sn_4_19 '0*vdd + 1*vss'
.DCVOLT sn_4_20 '0*vdd + 1*vss'
.DCVOLT sn_4_21 '0*vdd + 1*vss'
.DCVOLT sn_4_22 '0*vdd + 1*vss'
.DCVOLT sn_4_23 '0*vdd + 1*vss'
.DCVOLT sn_4_24 '0*vdd + 1*vss'
.DCVOLT sn_4_25 '0*vdd + 1*vss'
.DCVOLT sn_4_26 '0*vdd + 1*vss'
.DCVOLT sn_4_27 '0*vdd + 1*vss'
.DCVOLT sn_4_28 '0*vdd + 1*vss'
.DCVOLT sn_4_29 '0*vdd + 1*vss'
.DCVOLT sn_4_30 '0*vdd + 1*vss'
.DCVOLT sn_4_31 '0*vdd + 1*vss'
.DCVOLT sn_5_0 '0*vdd + 1*vss'
.DCVOLT sn_5_1 '0*vdd + 1*vss'
.DCVOLT sn_5_2 '0*vdd + 1*vss'
.DCVOLT sn_5_3 '0*vdd + 1*vss'
.DCVOLT sn_5_4 '0*vdd + 1*vss'
.DCVOLT sn_5_5 '0*vdd + 1*vss'
.DCVOLT sn_5_6 '0*vdd + 1*vss'
.DCVOLT sn_5_7 '0*vdd + 1*vss'
.DCVOLT sn_5_8 '0*vdd + 1*vss'
.DCVOLT sn_5_9 '0*vdd + 1*vss'
.DCVOLT sn_5_10 '0*vdd + 1*vss'
.DCVOLT sn_5_11 '0*vdd + 1*vss'
.DCVOLT sn_5_12 '0*vdd + 1*vss'
.DCVOLT sn_5_13 '0*vdd + 1*vss'
.DCVOLT sn_5_14 '0*vdd + 1*vss'
.DCVOLT sn_5_15 '0*vdd + 1*vss'
.DCVOLT sn_5_16 '0*vdd + 1*vss'
.DCVOLT sn_5_17 '0*vdd + 1*vss'
.DCVOLT sn_5_18 '0*vdd + 1*vss'
.DCVOLT sn_5_19 '0*vdd + 1*vss'
.DCVOLT sn_5_20 '0*vdd + 1*vss'
.DCVOLT sn_5_21 '0*vdd + 1*vss'
.DCVOLT sn_5_22 '0*vdd + 1*vss'
.DCVOLT sn_5_23 '0*vdd + 1*vss'
.DCVOLT sn_5_24 '0*vdd + 1*vss'
.DCVOLT sn_5_25 '0*vdd + 1*vss'
.DCVOLT sn_5_26 '0*vdd + 1*vss'
.DCVOLT sn_5_27 '0*vdd + 1*vss'
.DCVOLT sn_5_28 '0*vdd + 1*vss'
.DCVOLT sn_5_29 '0*vdd + 1*vss'
.DCVOLT sn_5_30 '0*vdd + 1*vss'
.DCVOLT sn_5_31 '0*vdd + 1*vss'
.DCVOLT sn_6_0 '0*vdd + 1*vss'
.DCVOLT sn_6_1 '0*vdd + 1*vss'
.DCVOLT sn_6_2 '0*vdd + 1*vss'
.DCVOLT sn_6_3 '0*vdd + 1*vss'
.DCVOLT sn_6_4 '0*vdd + 1*vss'
.DCVOLT sn_6_5 '0*vdd + 1*vss'
.DCVOLT sn_6_6 '0*vdd + 1*vss'
.DCVOLT sn_6_7 '0*vdd + 1*vss'
.DCVOLT sn_6_8 '0*vdd + 1*vss'
.DCVOLT sn_6_9 '0*vdd + 1*vss'
.DCVOLT sn_6_10 '0*vdd + 1*vss'
.DCVOLT sn_6_11 '0*vdd + 1*vss'
.DCVOLT sn_6_12 '0*vdd + 1*vss'
.DCVOLT sn_6_13 '0*vdd + 1*vss'
.DCVOLT sn_6_14 '0*vdd + 1*vss'
.DCVOLT sn_6_15 '0*vdd + 1*vss'
.DCVOLT sn_6_16 '0*vdd + 1*vss'
.DCVOLT sn_6_17 '0*vdd + 1*vss'
.DCVOLT sn_6_18 '0*vdd + 1*vss'
.DCVOLT sn_6_19 '0*vdd + 1*vss'
.DCVOLT sn_6_20 '0*vdd + 1*vss'
.DCVOLT sn_6_21 '0*vdd + 1*vss'
.DCVOLT sn_6_22 '0*vdd + 1*vss'
.DCVOLT sn_6_23 '0*vdd + 1*vss'
.DCVOLT sn_6_24 '0*vdd + 1*vss'
.DCVOLT sn_6_25 '0*vdd + 1*vss'
.DCVOLT sn_6_26 '0*vdd + 1*vss'
.DCVOLT sn_6_27 '0*vdd + 1*vss'
.DCVOLT sn_6_28 '0*vdd + 1*vss'
.DCVOLT sn_6_29 '0*vdd + 1*vss'
.DCVOLT sn_6_30 '0*vdd + 1*vss'
.DCVOLT sn_6_31 '0*vdd + 1*vss'
.DCVOLT sn_7_0 '0*vdd + 1*vss'
.DCVOLT sn_7_1 '0*vdd + 1*vss'
.DCVOLT sn_7_2 '0*vdd + 1*vss'
.DCVOLT sn_7_3 '0*vdd + 1*vss'
.DCVOLT sn_7_4 '0*vdd + 1*vss'
.DCVOLT sn_7_5 '0*vdd + 1*vss'
.DCVOLT sn_7_6 '0*vdd + 1*vss'
.DCVOLT sn_7_7 '0*vdd + 1*vss'
.DCVOLT sn_7_8 '0*vdd + 1*vss'
.DCVOLT sn_7_9 '0*vdd + 1*vss'
.DCVOLT sn_7_10 '0*vdd + 1*vss'
.DCVOLT sn_7_11 '0*vdd + 1*vss'
.DCVOLT sn_7_12 '0*vdd + 1*vss'
.DCVOLT sn_7_13 '0*vdd + 1*vss'
.DCVOLT sn_7_14 '0*vdd + 1*vss'
.DCVOLT sn_7_15 '0*vdd + 1*vss'
.DCVOLT sn_7_16 '0*vdd + 1*vss'
.DCVOLT sn_7_17 '0*vdd + 1*vss'
.DCVOLT sn_7_18 '0*vdd + 1*vss'
.DCVOLT sn_7_19 '0*vdd + 1*vss'
.DCVOLT sn_7_20 '0*vdd + 1*vss'
.DCVOLT sn_7_21 '0*vdd + 1*vss'
.DCVOLT sn_7_22 '0*vdd + 1*vss'
.DCVOLT sn_7_23 '0*vdd + 1*vss'
.DCVOLT sn_7_24 '0*vdd + 1*vss'
.DCVOLT sn_7_25 '0*vdd + 1*vss'
.DCVOLT sn_7_26 '0*vdd + 1*vss'
.DCVOLT sn_7_27 '0*vdd + 1*vss'
.DCVOLT sn_7_28 '0*vdd + 1*vss'
.DCVOLT sn_7_29 '0*vdd + 1*vss'
.DCVOLT sn_7_30 '0*vdd + 1*vss'
.DCVOLT sn_7_31 '0*vdd + 1*vss'
.DCVOLT sn_8_0 '0*vdd + 1*vss'
.DCVOLT sn_8_1 '0*vdd + 1*vss'
.DCVOLT sn_8_2 '0*vdd + 1*vss'
.DCVOLT sn_8_3 '0*vdd + 1*vss'
.DCVOLT sn_8_4 '0*vdd + 1*vss'
.DCVOLT sn_8_5 '0*vdd + 1*vss'
.DCVOLT sn_8_6 '0*vdd + 1*vss'
.DCVOLT sn_8_7 '0*vdd + 1*vss'
.DCVOLT sn_8_8 '0*vdd + 1*vss'
.DCVOLT sn_8_9 '0*vdd + 1*vss'
.DCVOLT sn_8_10 '0*vdd + 1*vss'
.DCVOLT sn_8_11 '0*vdd + 1*vss'
.DCVOLT sn_8_12 '0*vdd + 1*vss'
.DCVOLT sn_8_13 '0*vdd + 1*vss'
.DCVOLT sn_8_14 '0*vdd + 1*vss'
.DCVOLT sn_8_15 '0*vdd + 1*vss'
.DCVOLT sn_8_16 '0*vdd + 1*vss'
.DCVOLT sn_8_17 '0*vdd + 1*vss'
.DCVOLT sn_8_18 '0*vdd + 1*vss'
.DCVOLT sn_8_19 '0*vdd + 1*vss'
.DCVOLT sn_8_20 '0*vdd + 1*vss'
.DCVOLT sn_8_21 '0*vdd + 1*vss'
.DCVOLT sn_8_22 '0*vdd + 1*vss'
.DCVOLT sn_8_23 '0*vdd + 1*vss'
.DCVOLT sn_8_24 '0*vdd + 1*vss'
.DCVOLT sn_8_25 '0*vdd + 1*vss'
.DCVOLT sn_8_26 '0*vdd + 1*vss'
.DCVOLT sn_8_27 '0*vdd + 1*vss'
.DCVOLT sn_8_28 '0*vdd + 1*vss'
.DCVOLT sn_8_29 '0*vdd + 1*vss'
.DCVOLT sn_8_30 '0*vdd + 1*vss'
.DCVOLT sn_8_31 '0*vdd + 1*vss'
.DCVOLT sn_9_0 '0*vdd + 1*vss'
.DCVOLT sn_9_1 '0*vdd + 1*vss'
.DCVOLT sn_9_2 '0*vdd + 1*vss'
.DCVOLT sn_9_3 '0*vdd + 1*vss'
.DCVOLT sn_9_4 '0*vdd + 1*vss'
.DCVOLT sn_9_5 '0*vdd + 1*vss'
.DCVOLT sn_9_6 '0*vdd + 1*vss'
.DCVOLT sn_9_7 '0*vdd + 1*vss'
.DCVOLT sn_9_8 '0*vdd + 1*vss'
.DCVOLT sn_9_9 '0*vdd + 1*vss'
.DCVOLT sn_9_10 '0*vdd + 1*vss'
.DCVOLT sn_9_11 '0*vdd + 1*vss'
.DCVOLT sn_9_12 '0*vdd + 1*vss'
.DCVOLT sn_9_13 '0*vdd + 1*vss'
.DCVOLT sn_9_14 '0*vdd + 1*vss'
.DCVOLT sn_9_15 '0*vdd + 1*vss'
.DCVOLT sn_9_16 '0*vdd + 1*vss'
.DCVOLT sn_9_17 '0*vdd + 1*vss'
.DCVOLT sn_9_18 '0*vdd + 1*vss'
.DCVOLT sn_9_19 '0*vdd + 1*vss'
.DCVOLT sn_9_20 '0*vdd + 1*vss'
.DCVOLT sn_9_21 '0*vdd + 1*vss'
.DCVOLT sn_9_22 '0*vdd + 1*vss'
.DCVOLT sn_9_23 '0*vdd + 1*vss'
.DCVOLT sn_9_24 '0*vdd + 1*vss'
.DCVOLT sn_9_25 '0*vdd + 1*vss'
.DCVOLT sn_9_26 '0*vdd + 1*vss'
.DCVOLT sn_9_27 '0*vdd + 1*vss'
.DCVOLT sn_9_28 '0*vdd + 1*vss'
.DCVOLT sn_9_29 '0*vdd + 1*vss'
.DCVOLT sn_9_30 '0*vdd + 1*vss'
.DCVOLT sn_9_31 '0*vdd + 1*vss'
.DCVOLT sn_10_0 '0*vdd + 1*vss'
.DCVOLT sn_10_1 '0*vdd + 1*vss'
.DCVOLT sn_10_2 '0*vdd + 1*vss'
.DCVOLT sn_10_3 '0*vdd + 1*vss'
.DCVOLT sn_10_4 '0*vdd + 1*vss'
.DCVOLT sn_10_5 '0*vdd + 1*vss'
.DCVOLT sn_10_6 '0*vdd + 1*vss'
.DCVOLT sn_10_7 '0*vdd + 1*vss'
.DCVOLT sn_10_8 '0*vdd + 1*vss'
.DCVOLT sn_10_9 '0*vdd + 1*vss'
.DCVOLT sn_10_10 '0*vdd + 1*vss'
.DCVOLT sn_10_11 '0*vdd + 1*vss'
.DCVOLT sn_10_12 '0*vdd + 1*vss'
.DCVOLT sn_10_13 '0*vdd + 1*vss'
.DCVOLT sn_10_14 '0*vdd + 1*vss'
.DCVOLT sn_10_15 '0*vdd + 1*vss'
.DCVOLT sn_10_16 '0*vdd + 1*vss'
.DCVOLT sn_10_17 '0*vdd + 1*vss'
.DCVOLT sn_10_18 '0*vdd + 1*vss'
.DCVOLT sn_10_19 '0*vdd + 1*vss'
.DCVOLT sn_10_20 '0*vdd + 1*vss'
.DCVOLT sn_10_21 '0*vdd + 1*vss'
.DCVOLT sn_10_22 '0*vdd + 1*vss'
.DCVOLT sn_10_23 '0*vdd + 1*vss'
.DCVOLT sn_10_24 '0*vdd + 1*vss'
.DCVOLT sn_10_25 '0*vdd + 1*vss'
.DCVOLT sn_10_26 '0*vdd + 1*vss'
.DCVOLT sn_10_27 '0*vdd + 1*vss'
.DCVOLT sn_10_28 '0*vdd + 1*vss'
.DCVOLT sn_10_29 '0*vdd + 1*vss'
.DCVOLT sn_10_30 '0*vdd + 1*vss'
.DCVOLT sn_10_31 '0*vdd + 1*vss'
.DCVOLT sn_11_0 '0*vdd + 1*vss'
.DCVOLT sn_11_1 '0*vdd + 1*vss'
.DCVOLT sn_11_2 '0*vdd + 1*vss'
.DCVOLT sn_11_3 '0*vdd + 1*vss'
.DCVOLT sn_11_4 '0*vdd + 1*vss'
.DCVOLT sn_11_5 '0*vdd + 1*vss'
.DCVOLT sn_11_6 '0*vdd + 1*vss'
.DCVOLT sn_11_7 '0*vdd + 1*vss'
.DCVOLT sn_11_8 '0*vdd + 1*vss'
.DCVOLT sn_11_9 '0*vdd + 1*vss'
.DCVOLT sn_11_10 '0*vdd + 1*vss'
.DCVOLT sn_11_11 '0*vdd + 1*vss'
.DCVOLT sn_11_12 '0*vdd + 1*vss'
.DCVOLT sn_11_13 '0*vdd + 1*vss'
.DCVOLT sn_11_14 '0*vdd + 1*vss'
.DCVOLT sn_11_15 '0*vdd + 1*vss'
.DCVOLT sn_11_16 '0*vdd + 1*vss'
.DCVOLT sn_11_17 '0*vdd + 1*vss'
.DCVOLT sn_11_18 '0*vdd + 1*vss'
.DCVOLT sn_11_19 '0*vdd + 1*vss'
.DCVOLT sn_11_20 '0*vdd + 1*vss'
.DCVOLT sn_11_21 '0*vdd + 1*vss'
.DCVOLT sn_11_22 '0*vdd + 1*vss'
.DCVOLT sn_11_23 '0*vdd + 1*vss'
.DCVOLT sn_11_24 '0*vdd + 1*vss'
.DCVOLT sn_11_25 '0*vdd + 1*vss'
.DCVOLT sn_11_26 '0*vdd + 1*vss'
.DCVOLT sn_11_27 '0*vdd + 1*vss'
.DCVOLT sn_11_28 '0*vdd + 1*vss'
.DCVOLT sn_11_29 '0*vdd + 1*vss'
.DCVOLT sn_11_30 '0*vdd + 1*vss'
.DCVOLT sn_11_31 '0*vdd + 1*vss'
.DCVOLT sn_12_0 '0*vdd + 1*vss'
.DCVOLT sn_12_1 '0*vdd + 1*vss'
.DCVOLT sn_12_2 '0*vdd + 1*vss'
.DCVOLT sn_12_3 '0*vdd + 1*vss'
.DCVOLT sn_12_4 '0*vdd + 1*vss'
.DCVOLT sn_12_5 '0*vdd + 1*vss'
.DCVOLT sn_12_6 '0*vdd + 1*vss'
.DCVOLT sn_12_7 '0*vdd + 1*vss'
.DCVOLT sn_12_8 '0*vdd + 1*vss'
.DCVOLT sn_12_9 '0*vdd + 1*vss'
.DCVOLT sn_12_10 '0*vdd + 1*vss'
.DCVOLT sn_12_11 '0*vdd + 1*vss'
.DCVOLT sn_12_12 '0*vdd + 1*vss'
.DCVOLT sn_12_13 '0*vdd + 1*vss'
.DCVOLT sn_12_14 '0*vdd + 1*vss'
.DCVOLT sn_12_15 '0*vdd + 1*vss'
.DCVOLT sn_12_16 '0*vdd + 1*vss'
.DCVOLT sn_12_17 '0*vdd + 1*vss'
.DCVOLT sn_12_18 '0*vdd + 1*vss'
.DCVOLT sn_12_19 '0*vdd + 1*vss'
.DCVOLT sn_12_20 '0*vdd + 1*vss'
.DCVOLT sn_12_21 '0*vdd + 1*vss'
.DCVOLT sn_12_22 '0*vdd + 1*vss'
.DCVOLT sn_12_23 '0*vdd + 1*vss'
.DCVOLT sn_12_24 '0*vdd + 1*vss'
.DCVOLT sn_12_25 '0*vdd + 1*vss'
.DCVOLT sn_12_26 '0*vdd + 1*vss'
.DCVOLT sn_12_27 '0*vdd + 1*vss'
.DCVOLT sn_12_28 '0*vdd + 1*vss'
.DCVOLT sn_12_29 '0*vdd + 1*vss'
.DCVOLT sn_12_30 '0*vdd + 1*vss'
.DCVOLT sn_12_31 '0*vdd + 1*vss'
.DCVOLT sn_13_0 '0*vdd + 1*vss'
.DCVOLT sn_13_1 '0*vdd + 1*vss'
.DCVOLT sn_13_2 '0*vdd + 1*vss'
.DCVOLT sn_13_3 '0*vdd + 1*vss'
.DCVOLT sn_13_4 '0*vdd + 1*vss'
.DCVOLT sn_13_5 '0*vdd + 1*vss'
.DCVOLT sn_13_6 '0*vdd + 1*vss'
.DCVOLT sn_13_7 '0*vdd + 1*vss'
.DCVOLT sn_13_8 '0*vdd + 1*vss'
.DCVOLT sn_13_9 '0*vdd + 1*vss'
.DCVOLT sn_13_10 '0*vdd + 1*vss'
.DCVOLT sn_13_11 '0*vdd + 1*vss'
.DCVOLT sn_13_12 '0*vdd + 1*vss'
.DCVOLT sn_13_13 '0*vdd + 1*vss'
.DCVOLT sn_13_14 '0*vdd + 1*vss'
.DCVOLT sn_13_15 '0*vdd + 1*vss'
.DCVOLT sn_13_16 '0*vdd + 1*vss'
.DCVOLT sn_13_17 '0*vdd + 1*vss'
.DCVOLT sn_13_18 '0*vdd + 1*vss'
.DCVOLT sn_13_19 '0*vdd + 1*vss'
.DCVOLT sn_13_20 '0*vdd + 1*vss'
.DCVOLT sn_13_21 '0*vdd + 1*vss'
.DCVOLT sn_13_22 '0*vdd + 1*vss'
.DCVOLT sn_13_23 '0*vdd + 1*vss'
.DCVOLT sn_13_24 '0*vdd + 1*vss'
.DCVOLT sn_13_25 '0*vdd + 1*vss'
.DCVOLT sn_13_26 '0*vdd + 1*vss'
.DCVOLT sn_13_27 '0*vdd + 1*vss'
.DCVOLT sn_13_28 '0*vdd + 1*vss'
.DCVOLT sn_13_29 '0*vdd + 1*vss'
.DCVOLT sn_13_30 '0*vdd + 1*vss'
.DCVOLT sn_13_31 '0*vdd + 1*vss'
.DCVOLT sn_14_0 '0*vdd + 1*vss'
.DCVOLT sn_14_1 '0*vdd + 1*vss'
.DCVOLT sn_14_2 '0*vdd + 1*vss'
.DCVOLT sn_14_3 '0*vdd + 1*vss'
.DCVOLT sn_14_4 '0*vdd + 1*vss'
.DCVOLT sn_14_5 '0*vdd + 1*vss'
.DCVOLT sn_14_6 '0*vdd + 1*vss'
.DCVOLT sn_14_7 '0*vdd + 1*vss'
.DCVOLT sn_14_8 '0*vdd + 1*vss'
.DCVOLT sn_14_9 '0*vdd + 1*vss'
.DCVOLT sn_14_10 '0*vdd + 1*vss'
.DCVOLT sn_14_11 '0*vdd + 1*vss'
.DCVOLT sn_14_12 '0*vdd + 1*vss'
.DCVOLT sn_14_13 '0*vdd + 1*vss'
.DCVOLT sn_14_14 '0*vdd + 1*vss'
.DCVOLT sn_14_15 '0*vdd + 1*vss'
.DCVOLT sn_14_16 '0*vdd + 1*vss'
.DCVOLT sn_14_17 '0*vdd + 1*vss'
.DCVOLT sn_14_18 '0*vdd + 1*vss'
.DCVOLT sn_14_19 '0*vdd + 1*vss'
.DCVOLT sn_14_20 '0*vdd + 1*vss'
.DCVOLT sn_14_21 '0*vdd + 1*vss'
.DCVOLT sn_14_22 '0*vdd + 1*vss'
.DCVOLT sn_14_23 '0*vdd + 1*vss'
.DCVOLT sn_14_24 '0*vdd + 1*vss'
.DCVOLT sn_14_25 '0*vdd + 1*vss'
.DCVOLT sn_14_26 '0*vdd + 1*vss'
.DCVOLT sn_14_27 '0*vdd + 1*vss'
.DCVOLT sn_14_28 '0*vdd + 1*vss'
.DCVOLT sn_14_29 '0*vdd + 1*vss'
.DCVOLT sn_14_30 '0*vdd + 1*vss'
.DCVOLT sn_14_31 '0*vdd + 1*vss'
.DCVOLT sn_15_0 '0*vdd + 1*vss'
.DCVOLT sn_15_1 '0*vdd + 1*vss'
.DCVOLT sn_15_2 '0*vdd + 1*vss'
.DCVOLT sn_15_3 '0*vdd + 1*vss'
.DCVOLT sn_15_4 '0*vdd + 1*vss'
.DCVOLT sn_15_5 '0*vdd + 1*vss'
.DCVOLT sn_15_6 '0*vdd + 1*vss'
.DCVOLT sn_15_7 '0*vdd + 1*vss'
.DCVOLT sn_15_8 '0*vdd + 1*vss'
.DCVOLT sn_15_9 '0*vdd + 1*vss'
.DCVOLT sn_15_10 '0*vdd + 1*vss'
.DCVOLT sn_15_11 '0*vdd + 1*vss'
.DCVOLT sn_15_12 '0*vdd + 1*vss'
.DCVOLT sn_15_13 '0*vdd + 1*vss'
.DCVOLT sn_15_14 '0*vdd + 1*vss'
.DCVOLT sn_15_15 '0*vdd + 1*vss'
.DCVOLT sn_15_16 '0*vdd + 1*vss'
.DCVOLT sn_15_17 '0*vdd + 1*vss'
.DCVOLT sn_15_18 '0*vdd + 1*vss'
.DCVOLT sn_15_19 '0*vdd + 1*vss'
.DCVOLT sn_15_20 '0*vdd + 1*vss'
.DCVOLT sn_15_21 '0*vdd + 1*vss'
.DCVOLT sn_15_22 '0*vdd + 1*vss'
.DCVOLT sn_15_23 '0*vdd + 1*vss'
.DCVOLT sn_15_24 '0*vdd + 1*vss'
.DCVOLT sn_15_25 '0*vdd + 1*vss'
.DCVOLT sn_15_26 '0*vdd + 1*vss'
.DCVOLT sn_15_27 '0*vdd + 1*vss'
.DCVOLT sn_15_28 '0*vdd + 1*vss'
.DCVOLT sn_15_29 '0*vdd + 1*vss'
.DCVOLT sn_15_30 '0*vdd + 1*vss'
.DCVOLT sn_15_31 '0*vdd + 1*vss'
.DCVOLT sn_16_0 '0*vdd + 1*vss'
.DCVOLT sn_16_1 '0*vdd + 1*vss'
.DCVOLT sn_16_2 '0*vdd + 1*vss'
.DCVOLT sn_16_3 '0*vdd + 1*vss'
.DCVOLT sn_16_4 '0*vdd + 1*vss'
.DCVOLT sn_16_5 '0*vdd + 1*vss'
.DCVOLT sn_16_6 '0*vdd + 1*vss'
.DCVOLT sn_16_7 '0*vdd + 1*vss'
.DCVOLT sn_16_8 '0*vdd + 1*vss'
.DCVOLT sn_16_9 '0*vdd + 1*vss'
.DCVOLT sn_16_10 '0*vdd + 1*vss'
.DCVOLT sn_16_11 '0*vdd + 1*vss'
.DCVOLT sn_16_12 '0*vdd + 1*vss'
.DCVOLT sn_16_13 '0*vdd + 1*vss'
.DCVOLT sn_16_14 '0*vdd + 1*vss'
.DCVOLT sn_16_15 '0*vdd + 1*vss'
.DCVOLT sn_16_16 '0*vdd + 1*vss'
.DCVOLT sn_16_17 '0*vdd + 1*vss'
.DCVOLT sn_16_18 '0*vdd + 1*vss'
.DCVOLT sn_16_19 '0*vdd + 1*vss'
.DCVOLT sn_16_20 '0*vdd + 1*vss'
.DCVOLT sn_16_21 '0*vdd + 1*vss'
.DCVOLT sn_16_22 '0*vdd + 1*vss'
.DCVOLT sn_16_23 '0*vdd + 1*vss'
.DCVOLT sn_16_24 '0*vdd + 1*vss'
.DCVOLT sn_16_25 '0*vdd + 1*vss'
.DCVOLT sn_16_26 '0*vdd + 1*vss'
.DCVOLT sn_16_27 '0*vdd + 1*vss'
.DCVOLT sn_16_28 '0*vdd + 1*vss'
.DCVOLT sn_16_29 '0*vdd + 1*vss'
.DCVOLT sn_16_30 '0*vdd + 1*vss'
.DCVOLT sn_16_31 '0*vdd + 1*vss'
.DCVOLT sn_17_0 '0*vdd + 1*vss'
.DCVOLT sn_17_1 '0*vdd + 1*vss'
.DCVOLT sn_17_2 '0*vdd + 1*vss'
.DCVOLT sn_17_3 '0*vdd + 1*vss'
.DCVOLT sn_17_4 '0*vdd + 1*vss'
.DCVOLT sn_17_5 '0*vdd + 1*vss'
.DCVOLT sn_17_6 '0*vdd + 1*vss'
.DCVOLT sn_17_7 '0*vdd + 1*vss'
.DCVOLT sn_17_8 '0*vdd + 1*vss'
.DCVOLT sn_17_9 '0*vdd + 1*vss'
.DCVOLT sn_17_10 '0*vdd + 1*vss'
.DCVOLT sn_17_11 '0*vdd + 1*vss'
.DCVOLT sn_17_12 '0*vdd + 1*vss'
.DCVOLT sn_17_13 '0*vdd + 1*vss'
.DCVOLT sn_17_14 '0*vdd + 1*vss'
.DCVOLT sn_17_15 '0*vdd + 1*vss'
.DCVOLT sn_17_16 '0*vdd + 1*vss'
.DCVOLT sn_17_17 '0*vdd + 1*vss'
.DCVOLT sn_17_18 '0*vdd + 1*vss'
.DCVOLT sn_17_19 '0*vdd + 1*vss'
.DCVOLT sn_17_20 '0*vdd + 1*vss'
.DCVOLT sn_17_21 '0*vdd + 1*vss'
.DCVOLT sn_17_22 '0*vdd + 1*vss'
.DCVOLT sn_17_23 '0*vdd + 1*vss'
.DCVOLT sn_17_24 '0*vdd + 1*vss'
.DCVOLT sn_17_25 '0*vdd + 1*vss'
.DCVOLT sn_17_26 '0*vdd + 1*vss'
.DCVOLT sn_17_27 '0*vdd + 1*vss'
.DCVOLT sn_17_28 '0*vdd + 1*vss'
.DCVOLT sn_17_29 '0*vdd + 1*vss'
.DCVOLT sn_17_30 '0*vdd + 1*vss'
.DCVOLT sn_17_31 '0*vdd + 1*vss'
.DCVOLT sn_18_0 '0*vdd + 1*vss'
.DCVOLT sn_18_1 '0*vdd + 1*vss'
.DCVOLT sn_18_2 '0*vdd + 1*vss'
.DCVOLT sn_18_3 '0*vdd + 1*vss'
.DCVOLT sn_18_4 '0*vdd + 1*vss'
.DCVOLT sn_18_5 '0*vdd + 1*vss'
.DCVOLT sn_18_6 '0*vdd + 1*vss'
.DCVOLT sn_18_7 '0*vdd + 1*vss'
.DCVOLT sn_18_8 '0*vdd + 1*vss'
.DCVOLT sn_18_9 '0*vdd + 1*vss'
.DCVOLT sn_18_10 '0*vdd + 1*vss'
.DCVOLT sn_18_11 '0*vdd + 1*vss'
.DCVOLT sn_18_12 '0*vdd + 1*vss'
.DCVOLT sn_18_13 '0*vdd + 1*vss'
.DCVOLT sn_18_14 '0*vdd + 1*vss'
.DCVOLT sn_18_15 '0*vdd + 1*vss'
.DCVOLT sn_18_16 '0*vdd + 1*vss'
.DCVOLT sn_18_17 '0*vdd + 1*vss'
.DCVOLT sn_18_18 '0*vdd + 1*vss'
.DCVOLT sn_18_19 '0*vdd + 1*vss'
.DCVOLT sn_18_20 '0*vdd + 1*vss'
.DCVOLT sn_18_21 '0*vdd + 1*vss'
.DCVOLT sn_18_22 '0*vdd + 1*vss'
.DCVOLT sn_18_23 '0*vdd + 1*vss'
.DCVOLT sn_18_24 '0*vdd + 1*vss'
.DCVOLT sn_18_25 '0*vdd + 1*vss'
.DCVOLT sn_18_26 '0*vdd + 1*vss'
.DCVOLT sn_18_27 '0*vdd + 1*vss'
.DCVOLT sn_18_28 '0*vdd + 1*vss'
.DCVOLT sn_18_29 '0*vdd + 1*vss'
.DCVOLT sn_18_30 '0*vdd + 1*vss'
.DCVOLT sn_18_31 '0*vdd + 1*vss'
.DCVOLT sn_19_0 '0*vdd + 1*vss'
.DCVOLT sn_19_1 '0*vdd + 1*vss'
.DCVOLT sn_19_2 '0*vdd + 1*vss'
.DCVOLT sn_19_3 '0*vdd + 1*vss'
.DCVOLT sn_19_4 '0*vdd + 1*vss'
.DCVOLT sn_19_5 '0*vdd + 1*vss'
.DCVOLT sn_19_6 '0*vdd + 1*vss'
.DCVOLT sn_19_7 '0*vdd + 1*vss'
.DCVOLT sn_19_8 '0*vdd + 1*vss'
.DCVOLT sn_19_9 '0*vdd + 1*vss'
.DCVOLT sn_19_10 '0*vdd + 1*vss'
.DCVOLT sn_19_11 '0*vdd + 1*vss'
.DCVOLT sn_19_12 '0*vdd + 1*vss'
.DCVOLT sn_19_13 '0*vdd + 1*vss'
.DCVOLT sn_19_14 '0*vdd + 1*vss'
.DCVOLT sn_19_15 '0*vdd + 1*vss'
.DCVOLT sn_19_16 '0*vdd + 1*vss'
.DCVOLT sn_19_17 '0*vdd + 1*vss'
.DCVOLT sn_19_18 '0*vdd + 1*vss'
.DCVOLT sn_19_19 '0*vdd + 1*vss'
.DCVOLT sn_19_20 '0*vdd + 1*vss'
.DCVOLT sn_19_21 '0*vdd + 1*vss'
.DCVOLT sn_19_22 '0*vdd + 1*vss'
.DCVOLT sn_19_23 '0*vdd + 1*vss'
.DCVOLT sn_19_24 '0*vdd + 1*vss'
.DCVOLT sn_19_25 '0*vdd + 1*vss'
.DCVOLT sn_19_26 '0*vdd + 1*vss'
.DCVOLT sn_19_27 '0*vdd + 1*vss'
.DCVOLT sn_19_28 '0*vdd + 1*vss'
.DCVOLT sn_19_29 '0*vdd + 1*vss'
.DCVOLT sn_19_30 '0*vdd + 1*vss'
.DCVOLT sn_19_31 '0*vdd + 1*vss'
.DCVOLT sn_20_0 '0*vdd + 1*vss'
.DCVOLT sn_20_1 '0*vdd + 1*vss'
.DCVOLT sn_20_2 '0*vdd + 1*vss'
.DCVOLT sn_20_3 '0*vdd + 1*vss'
.DCVOLT sn_20_4 '0*vdd + 1*vss'
.DCVOLT sn_20_5 '0*vdd + 1*vss'
.DCVOLT sn_20_6 '0*vdd + 1*vss'
.DCVOLT sn_20_7 '0*vdd + 1*vss'
.DCVOLT sn_20_8 '0*vdd + 1*vss'
.DCVOLT sn_20_9 '0*vdd + 1*vss'
.DCVOLT sn_20_10 '0*vdd + 1*vss'
.DCVOLT sn_20_11 '0*vdd + 1*vss'
.DCVOLT sn_20_12 '0*vdd + 1*vss'
.DCVOLT sn_20_13 '0*vdd + 1*vss'
.DCVOLT sn_20_14 '0*vdd + 1*vss'
.DCVOLT sn_20_15 '0*vdd + 1*vss'
.DCVOLT sn_20_16 '0*vdd + 1*vss'
.DCVOLT sn_20_17 '0*vdd + 1*vss'
.DCVOLT sn_20_18 '0*vdd + 1*vss'
.DCVOLT sn_20_19 '0*vdd + 1*vss'
.DCVOLT sn_20_20 '0*vdd + 1*vss'
.DCVOLT sn_20_21 '0*vdd + 1*vss'
.DCVOLT sn_20_22 '0*vdd + 1*vss'
.DCVOLT sn_20_23 '0*vdd + 1*vss'
.DCVOLT sn_20_24 '0*vdd + 1*vss'
.DCVOLT sn_20_25 '0*vdd + 1*vss'
.DCVOLT sn_20_26 '0*vdd + 1*vss'
.DCVOLT sn_20_27 '0*vdd + 1*vss'
.DCVOLT sn_20_28 '0*vdd + 1*vss'
.DCVOLT sn_20_29 '0*vdd + 1*vss'
.DCVOLT sn_20_30 '0*vdd + 1*vss'
.DCVOLT sn_20_31 '0*vdd + 1*vss'
.DCVOLT sn_21_0 '0*vdd + 1*vss'
.DCVOLT sn_21_1 '0*vdd + 1*vss'
.DCVOLT sn_21_2 '0*vdd + 1*vss'
.DCVOLT sn_21_3 '0*vdd + 1*vss'
.DCVOLT sn_21_4 '0*vdd + 1*vss'
.DCVOLT sn_21_5 '0*vdd + 1*vss'
.DCVOLT sn_21_6 '0*vdd + 1*vss'
.DCVOLT sn_21_7 '0*vdd + 1*vss'
.DCVOLT sn_21_8 '0*vdd + 1*vss'
.DCVOLT sn_21_9 '0*vdd + 1*vss'
.DCVOLT sn_21_10 '0*vdd + 1*vss'
.DCVOLT sn_21_11 '0*vdd + 1*vss'
.DCVOLT sn_21_12 '0*vdd + 1*vss'
.DCVOLT sn_21_13 '0*vdd + 1*vss'
.DCVOLT sn_21_14 '0*vdd + 1*vss'
.DCVOLT sn_21_15 '0*vdd + 1*vss'
.DCVOLT sn_21_16 '0*vdd + 1*vss'
.DCVOLT sn_21_17 '0*vdd + 1*vss'
.DCVOLT sn_21_18 '0*vdd + 1*vss'
.DCVOLT sn_21_19 '0*vdd + 1*vss'
.DCVOLT sn_21_20 '0*vdd + 1*vss'
.DCVOLT sn_21_21 '0*vdd + 1*vss'
.DCVOLT sn_21_22 '0*vdd + 1*vss'
.DCVOLT sn_21_23 '0*vdd + 1*vss'
.DCVOLT sn_21_24 '0*vdd + 1*vss'
.DCVOLT sn_21_25 '0*vdd + 1*vss'
.DCVOLT sn_21_26 '0*vdd + 1*vss'
.DCVOLT sn_21_27 '0*vdd + 1*vss'
.DCVOLT sn_21_28 '0*vdd + 1*vss'
.DCVOLT sn_21_29 '0*vdd + 1*vss'
.DCVOLT sn_21_30 '0*vdd + 1*vss'
.DCVOLT sn_21_31 '0*vdd + 1*vss'
.DCVOLT sn_22_0 '0*vdd + 1*vss'
.DCVOLT sn_22_1 '0*vdd + 1*vss'
.DCVOLT sn_22_2 '0*vdd + 1*vss'
.DCVOLT sn_22_3 '0*vdd + 1*vss'
.DCVOLT sn_22_4 '0*vdd + 1*vss'
.DCVOLT sn_22_5 '0*vdd + 1*vss'
.DCVOLT sn_22_6 '0*vdd + 1*vss'
.DCVOLT sn_22_7 '0*vdd + 1*vss'
.DCVOLT sn_22_8 '0*vdd + 1*vss'
.DCVOLT sn_22_9 '0*vdd + 1*vss'
.DCVOLT sn_22_10 '0*vdd + 1*vss'
.DCVOLT sn_22_11 '0*vdd + 1*vss'
.DCVOLT sn_22_12 '0*vdd + 1*vss'
.DCVOLT sn_22_13 '0*vdd + 1*vss'
.DCVOLT sn_22_14 '0*vdd + 1*vss'
.DCVOLT sn_22_15 '0*vdd + 1*vss'
.DCVOLT sn_22_16 '0*vdd + 1*vss'
.DCVOLT sn_22_17 '0*vdd + 1*vss'
.DCVOLT sn_22_18 '0*vdd + 1*vss'
.DCVOLT sn_22_19 '0*vdd + 1*vss'
.DCVOLT sn_22_20 '0*vdd + 1*vss'
.DCVOLT sn_22_21 '0*vdd + 1*vss'
.DCVOLT sn_22_22 '0*vdd + 1*vss'
.DCVOLT sn_22_23 '0*vdd + 1*vss'
.DCVOLT sn_22_24 '0*vdd + 1*vss'
.DCVOLT sn_22_25 '0*vdd + 1*vss'
.DCVOLT sn_22_26 '0*vdd + 1*vss'
.DCVOLT sn_22_27 '0*vdd + 1*vss'
.DCVOLT sn_22_28 '0*vdd + 1*vss'
.DCVOLT sn_22_29 '0*vdd + 1*vss'
.DCVOLT sn_22_30 '0*vdd + 1*vss'
.DCVOLT sn_22_31 '0*vdd + 1*vss'
.DCVOLT sn_23_0 '0*vdd + 1*vss'
.DCVOLT sn_23_1 '0*vdd + 1*vss'
.DCVOLT sn_23_2 '0*vdd + 1*vss'
.DCVOLT sn_23_3 '0*vdd + 1*vss'
.DCVOLT sn_23_4 '0*vdd + 1*vss'
.DCVOLT sn_23_5 '0*vdd + 1*vss'
.DCVOLT sn_23_6 '0*vdd + 1*vss'
.DCVOLT sn_23_7 '0*vdd + 1*vss'
.DCVOLT sn_23_8 '0*vdd + 1*vss'
.DCVOLT sn_23_9 '0*vdd + 1*vss'
.DCVOLT sn_23_10 '0*vdd + 1*vss'
.DCVOLT sn_23_11 '0*vdd + 1*vss'
.DCVOLT sn_23_12 '0*vdd + 1*vss'
.DCVOLT sn_23_13 '0*vdd + 1*vss'
.DCVOLT sn_23_14 '0*vdd + 1*vss'
.DCVOLT sn_23_15 '0*vdd + 1*vss'
.DCVOLT sn_23_16 '0*vdd + 1*vss'
.DCVOLT sn_23_17 '0*vdd + 1*vss'
.DCVOLT sn_23_18 '0*vdd + 1*vss'
.DCVOLT sn_23_19 '0*vdd + 1*vss'
.DCVOLT sn_23_20 '0*vdd + 1*vss'
.DCVOLT sn_23_21 '0*vdd + 1*vss'
.DCVOLT sn_23_22 '0*vdd + 1*vss'
.DCVOLT sn_23_23 '0*vdd + 1*vss'
.DCVOLT sn_23_24 '0*vdd + 1*vss'
.DCVOLT sn_23_25 '0*vdd + 1*vss'
.DCVOLT sn_23_26 '0*vdd + 1*vss'
.DCVOLT sn_23_27 '0*vdd + 1*vss'
.DCVOLT sn_23_28 '0*vdd + 1*vss'
.DCVOLT sn_23_29 '0*vdd + 1*vss'
.DCVOLT sn_23_30 '0*vdd + 1*vss'
.DCVOLT sn_23_31 '0*vdd + 1*vss'
.DCVOLT sn_24_0 '0*vdd + 1*vss'
.DCVOLT sn_24_1 '0*vdd + 1*vss'
.DCVOLT sn_24_2 '0*vdd + 1*vss'
.DCVOLT sn_24_3 '0*vdd + 1*vss'
.DCVOLT sn_24_4 '0*vdd + 1*vss'
.DCVOLT sn_24_5 '0*vdd + 1*vss'
.DCVOLT sn_24_6 '0*vdd + 1*vss'
.DCVOLT sn_24_7 '0*vdd + 1*vss'
.DCVOLT sn_24_8 '0*vdd + 1*vss'
.DCVOLT sn_24_9 '0*vdd + 1*vss'
.DCVOLT sn_24_10 '0*vdd + 1*vss'
.DCVOLT sn_24_11 '0*vdd + 1*vss'
.DCVOLT sn_24_12 '0*vdd + 1*vss'
.DCVOLT sn_24_13 '0*vdd + 1*vss'
.DCVOLT sn_24_14 '0*vdd + 1*vss'
.DCVOLT sn_24_15 '0*vdd + 1*vss'
.DCVOLT sn_24_16 '0*vdd + 1*vss'
.DCVOLT sn_24_17 '0*vdd + 1*vss'
.DCVOLT sn_24_18 '0*vdd + 1*vss'
.DCVOLT sn_24_19 '0*vdd + 1*vss'
.DCVOLT sn_24_20 '0*vdd + 1*vss'
.DCVOLT sn_24_21 '0*vdd + 1*vss'
.DCVOLT sn_24_22 '0*vdd + 1*vss'
.DCVOLT sn_24_23 '0*vdd + 1*vss'
.DCVOLT sn_24_24 '0*vdd + 1*vss'
.DCVOLT sn_24_25 '0*vdd + 1*vss'
.DCVOLT sn_24_26 '0*vdd + 1*vss'
.DCVOLT sn_24_27 '0*vdd + 1*vss'
.DCVOLT sn_24_28 '0*vdd + 1*vss'
.DCVOLT sn_24_29 '0*vdd + 1*vss'
.DCVOLT sn_24_30 '0*vdd + 1*vss'
.DCVOLT sn_24_31 '0*vdd + 1*vss'
.DCVOLT sn_25_0 '0*vdd + 1*vss'
.DCVOLT sn_25_1 '0*vdd + 1*vss'
.DCVOLT sn_25_2 '0*vdd + 1*vss'
.DCVOLT sn_25_3 '0*vdd + 1*vss'
.DCVOLT sn_25_4 '0*vdd + 1*vss'
.DCVOLT sn_25_5 '0*vdd + 1*vss'
.DCVOLT sn_25_6 '0*vdd + 1*vss'
.DCVOLT sn_25_7 '0*vdd + 1*vss'
.DCVOLT sn_25_8 '0*vdd + 1*vss'
.DCVOLT sn_25_9 '0*vdd + 1*vss'
.DCVOLT sn_25_10 '0*vdd + 1*vss'
.DCVOLT sn_25_11 '0*vdd + 1*vss'
.DCVOLT sn_25_12 '0*vdd + 1*vss'
.DCVOLT sn_25_13 '0*vdd + 1*vss'
.DCVOLT sn_25_14 '0*vdd + 1*vss'
.DCVOLT sn_25_15 '0*vdd + 1*vss'
.DCVOLT sn_25_16 '0*vdd + 1*vss'
.DCVOLT sn_25_17 '0*vdd + 1*vss'
.DCVOLT sn_25_18 '0*vdd + 1*vss'
.DCVOLT sn_25_19 '0*vdd + 1*vss'
.DCVOLT sn_25_20 '0*vdd + 1*vss'
.DCVOLT sn_25_21 '0*vdd + 1*vss'
.DCVOLT sn_25_22 '0*vdd + 1*vss'
.DCVOLT sn_25_23 '0*vdd + 1*vss'
.DCVOLT sn_25_24 '0*vdd + 1*vss'
.DCVOLT sn_25_25 '0*vdd + 1*vss'
.DCVOLT sn_25_26 '0*vdd + 1*vss'
.DCVOLT sn_25_27 '0*vdd + 1*vss'
.DCVOLT sn_25_28 '0*vdd + 1*vss'
.DCVOLT sn_25_29 '0*vdd + 1*vss'
.DCVOLT sn_25_30 '0*vdd + 1*vss'
.DCVOLT sn_25_31 '0*vdd + 1*vss'
.DCVOLT sn_26_0 '0*vdd + 1*vss'
.DCVOLT sn_26_1 '0*vdd + 1*vss'
.DCVOLT sn_26_2 '0*vdd + 1*vss'
.DCVOLT sn_26_3 '0*vdd + 1*vss'
.DCVOLT sn_26_4 '0*vdd + 1*vss'
.DCVOLT sn_26_5 '0*vdd + 1*vss'
.DCVOLT sn_26_6 '0*vdd + 1*vss'
.DCVOLT sn_26_7 '0*vdd + 1*vss'
.DCVOLT sn_26_8 '0*vdd + 1*vss'
.DCVOLT sn_26_9 '0*vdd + 1*vss'
.DCVOLT sn_26_10 '0*vdd + 1*vss'
.DCVOLT sn_26_11 '0*vdd + 1*vss'
.DCVOLT sn_26_12 '0*vdd + 1*vss'
.DCVOLT sn_26_13 '0*vdd + 1*vss'
.DCVOLT sn_26_14 '0*vdd + 1*vss'
.DCVOLT sn_26_15 '0*vdd + 1*vss'
.DCVOLT sn_26_16 '0*vdd + 1*vss'
.DCVOLT sn_26_17 '0*vdd + 1*vss'
.DCVOLT sn_26_18 '0*vdd + 1*vss'
.DCVOLT sn_26_19 '0*vdd + 1*vss'
.DCVOLT sn_26_20 '0*vdd + 1*vss'
.DCVOLT sn_26_21 '0*vdd + 1*vss'
.DCVOLT sn_26_22 '0*vdd + 1*vss'
.DCVOLT sn_26_23 '0*vdd + 1*vss'
.DCVOLT sn_26_24 '0*vdd + 1*vss'
.DCVOLT sn_26_25 '0*vdd + 1*vss'
.DCVOLT sn_26_26 '0*vdd + 1*vss'
.DCVOLT sn_26_27 '0*vdd + 1*vss'
.DCVOLT sn_26_28 '0*vdd + 1*vss'
.DCVOLT sn_26_29 '0*vdd + 1*vss'
.DCVOLT sn_26_30 '0*vdd + 1*vss'
.DCVOLT sn_26_31 '0*vdd + 1*vss'
.DCVOLT sn_27_0 '0*vdd + 1*vss'
.DCVOLT sn_27_1 '0*vdd + 1*vss'
.DCVOLT sn_27_2 '0*vdd + 1*vss'
.DCVOLT sn_27_3 '0*vdd + 1*vss'
.DCVOLT sn_27_4 '0*vdd + 1*vss'
.DCVOLT sn_27_5 '0*vdd + 1*vss'
.DCVOLT sn_27_6 '0*vdd + 1*vss'
.DCVOLT sn_27_7 '0*vdd + 1*vss'
.DCVOLT sn_27_8 '0*vdd + 1*vss'
.DCVOLT sn_27_9 '0*vdd + 1*vss'
.DCVOLT sn_27_10 '0*vdd + 1*vss'
.DCVOLT sn_27_11 '0*vdd + 1*vss'
.DCVOLT sn_27_12 '0*vdd + 1*vss'
.DCVOLT sn_27_13 '0*vdd + 1*vss'
.DCVOLT sn_27_14 '0*vdd + 1*vss'
.DCVOLT sn_27_15 '0*vdd + 1*vss'
.DCVOLT sn_27_16 '0*vdd + 1*vss'
.DCVOLT sn_27_17 '0*vdd + 1*vss'
.DCVOLT sn_27_18 '0*vdd + 1*vss'
.DCVOLT sn_27_19 '0*vdd + 1*vss'
.DCVOLT sn_27_20 '0*vdd + 1*vss'
.DCVOLT sn_27_21 '0*vdd + 1*vss'
.DCVOLT sn_27_22 '0*vdd + 1*vss'
.DCVOLT sn_27_23 '0*vdd + 1*vss'
.DCVOLT sn_27_24 '0*vdd + 1*vss'
.DCVOLT sn_27_25 '0*vdd + 1*vss'
.DCVOLT sn_27_26 '0*vdd + 1*vss'
.DCVOLT sn_27_27 '0*vdd + 1*vss'
.DCVOLT sn_27_28 '0*vdd + 1*vss'
.DCVOLT sn_27_29 '0*vdd + 1*vss'
.DCVOLT sn_27_30 '0*vdd + 1*vss'
.DCVOLT sn_27_31 '0*vdd + 1*vss'
.DCVOLT sn_28_0 '0*vdd + 1*vss'
.DCVOLT sn_28_1 '0*vdd + 1*vss'
.DCVOLT sn_28_2 '0*vdd + 1*vss'
.DCVOLT sn_28_3 '0*vdd + 1*vss'
.DCVOLT sn_28_4 '0*vdd + 1*vss'
.DCVOLT sn_28_5 '0*vdd + 1*vss'
.DCVOLT sn_28_6 '0*vdd + 1*vss'
.DCVOLT sn_28_7 '0*vdd + 1*vss'
.DCVOLT sn_28_8 '0*vdd + 1*vss'
.DCVOLT sn_28_9 '0*vdd + 1*vss'
.DCVOLT sn_28_10 '0*vdd + 1*vss'
.DCVOLT sn_28_11 '0*vdd + 1*vss'
.DCVOLT sn_28_12 '0*vdd + 1*vss'
.DCVOLT sn_28_13 '0*vdd + 1*vss'
.DCVOLT sn_28_14 '0*vdd + 1*vss'
.DCVOLT sn_28_15 '0*vdd + 1*vss'
.DCVOLT sn_28_16 '0*vdd + 1*vss'
.DCVOLT sn_28_17 '0*vdd + 1*vss'
.DCVOLT sn_28_18 '0*vdd + 1*vss'
.DCVOLT sn_28_19 '0*vdd + 1*vss'
.DCVOLT sn_28_20 '0*vdd + 1*vss'
.DCVOLT sn_28_21 '0*vdd + 1*vss'
.DCVOLT sn_28_22 '0*vdd + 1*vss'
.DCVOLT sn_28_23 '0*vdd + 1*vss'
.DCVOLT sn_28_24 '0*vdd + 1*vss'
.DCVOLT sn_28_25 '0*vdd + 1*vss'
.DCVOLT sn_28_26 '0*vdd + 1*vss'
.DCVOLT sn_28_27 '0*vdd + 1*vss'
.DCVOLT sn_28_28 '0*vdd + 1*vss'
.DCVOLT sn_28_29 '0*vdd + 1*vss'
.DCVOLT sn_28_30 '0*vdd + 1*vss'
.DCVOLT sn_28_31 '0*vdd + 1*vss'
.DCVOLT sn_29_0 '0*vdd + 1*vss'
.DCVOLT sn_29_1 '0*vdd + 1*vss'
.DCVOLT sn_29_2 '0*vdd + 1*vss'
.DCVOLT sn_29_3 '0*vdd + 1*vss'
.DCVOLT sn_29_4 '0*vdd + 1*vss'
.DCVOLT sn_29_5 '0*vdd + 1*vss'
.DCVOLT sn_29_6 '0*vdd + 1*vss'
.DCVOLT sn_29_7 '0*vdd + 1*vss'
.DCVOLT sn_29_8 '0*vdd + 1*vss'
.DCVOLT sn_29_9 '0*vdd + 1*vss'
.DCVOLT sn_29_10 '0*vdd + 1*vss'
.DCVOLT sn_29_11 '0*vdd + 1*vss'
.DCVOLT sn_29_12 '0*vdd + 1*vss'
.DCVOLT sn_29_13 '0*vdd + 1*vss'
.DCVOLT sn_29_14 '0*vdd + 1*vss'
.DCVOLT sn_29_15 '0*vdd + 1*vss'
.DCVOLT sn_29_16 '0*vdd + 1*vss'
.DCVOLT sn_29_17 '0*vdd + 1*vss'
.DCVOLT sn_29_18 '0*vdd + 1*vss'
.DCVOLT sn_29_19 '0*vdd + 1*vss'
.DCVOLT sn_29_20 '0*vdd + 1*vss'
.DCVOLT sn_29_21 '0*vdd + 1*vss'
.DCVOLT sn_29_22 '0*vdd + 1*vss'
.DCVOLT sn_29_23 '0*vdd + 1*vss'
.DCVOLT sn_29_24 '0*vdd + 1*vss'
.DCVOLT sn_29_25 '0*vdd + 1*vss'
.DCVOLT sn_29_26 '0*vdd + 1*vss'
.DCVOLT sn_29_27 '0*vdd + 1*vss'
.DCVOLT sn_29_28 '0*vdd + 1*vss'
.DCVOLT sn_29_29 '0*vdd + 1*vss'
.DCVOLT sn_29_30 '0*vdd + 1*vss'
.DCVOLT sn_29_31 '0*vdd + 1*vss'
.DCVOLT sn_30_0 '0*vdd + 1*vss'
.DCVOLT sn_30_1 '0*vdd + 1*vss'
.DCVOLT sn_30_2 '0*vdd + 1*vss'
.DCVOLT sn_30_3 '0*vdd + 1*vss'
.DCVOLT sn_30_4 '0*vdd + 1*vss'
.DCVOLT sn_30_5 '0*vdd + 1*vss'
.DCVOLT sn_30_6 '0*vdd + 1*vss'
.DCVOLT sn_30_7 '0*vdd + 1*vss'
.DCVOLT sn_30_8 '0*vdd + 1*vss'
.DCVOLT sn_30_9 '0*vdd + 1*vss'
.DCVOLT sn_30_10 '0*vdd + 1*vss'
.DCVOLT sn_30_11 '0*vdd + 1*vss'
.DCVOLT sn_30_12 '0*vdd + 1*vss'
.DCVOLT sn_30_13 '0*vdd + 1*vss'
.DCVOLT sn_30_14 '0*vdd + 1*vss'
.DCVOLT sn_30_15 '0*vdd + 1*vss'
.DCVOLT sn_30_16 '0*vdd + 1*vss'
.DCVOLT sn_30_17 '0*vdd + 1*vss'
.DCVOLT sn_30_18 '0*vdd + 1*vss'
.DCVOLT sn_30_19 '0*vdd + 1*vss'
.DCVOLT sn_30_20 '0*vdd + 1*vss'
.DCVOLT sn_30_21 '0*vdd + 1*vss'
.DCVOLT sn_30_22 '0*vdd + 1*vss'
.DCVOLT sn_30_23 '0*vdd + 1*vss'
.DCVOLT sn_30_24 '0*vdd + 1*vss'
.DCVOLT sn_30_25 '0*vdd + 1*vss'
.DCVOLT sn_30_26 '0*vdd + 1*vss'
.DCVOLT sn_30_27 '0*vdd + 1*vss'
.DCVOLT sn_30_28 '0*vdd + 1*vss'
.DCVOLT sn_30_29 '0*vdd + 1*vss'
.DCVOLT sn_30_30 '0*vdd + 1*vss'
.DCVOLT sn_30_31 '0*vdd + 1*vss'
.DCVOLT sn_31_0 '0*vdd + 1*vss'
.DCVOLT sn_31_1 '0*vdd + 1*vss'
.DCVOLT sn_31_2 '0*vdd + 1*vss'
.DCVOLT sn_31_3 '0*vdd + 1*vss'
.DCVOLT sn_31_4 '0*vdd + 1*vss'
.DCVOLT sn_31_5 '0*vdd + 1*vss'
.DCVOLT sn_31_6 '0*vdd + 1*vss'
.DCVOLT sn_31_7 '0*vdd + 1*vss'
.DCVOLT sn_31_8 '0*vdd + 1*vss'
.DCVOLT sn_31_9 '0*vdd + 1*vss'
.DCVOLT sn_31_10 '0*vdd + 1*vss'
.DCVOLT sn_31_11 '0*vdd + 1*vss'
.DCVOLT sn_31_12 '0*vdd + 1*vss'
.DCVOLT sn_31_13 '0*vdd + 1*vss'
.DCVOLT sn_31_14 '0*vdd + 1*vss'
.DCVOLT sn_31_15 '0*vdd + 1*vss'
.DCVOLT sn_31_16 '0*vdd + 1*vss'
.DCVOLT sn_31_17 '0*vdd + 1*vss'
.DCVOLT sn_31_18 '0*vdd + 1*vss'
.DCVOLT sn_31_19 '0*vdd + 1*vss'
.DCVOLT sn_31_20 '0*vdd + 1*vss'
.DCVOLT sn_31_21 '0*vdd + 1*vss'
.DCVOLT sn_31_22 '0*vdd + 1*vss'
.DCVOLT sn_31_23 '0*vdd + 1*vss'
.DCVOLT sn_31_24 '0*vdd + 1*vss'
.DCVOLT sn_31_25 '0*vdd + 1*vss'
.DCVOLT sn_31_26 '0*vdd + 1*vss'
.DCVOLT sn_31_27 '0*vdd + 1*vss'
.DCVOLT sn_31_28 '0*vdd + 1*vss'
.DCVOLT sn_31_29 '0*vdd + 1*vss'
.DCVOLT sn_31_30 '0*vdd + 1*vss'
.DCVOLT sn_31_31 '0*vdd + 1*vss'
xgc_0_0 wwl_0_0 wbl_0_0 rwl_0_0 rbl_0_0 sn_0_0 wos_ros_gc
xrc_wwl_0_0 wwl_0 wwl_0_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_0 wbl_0 wbl_0_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_0 rwl_0 rwl_0_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_0 rbl_0 rbl_0_0 rc_unit R0=Rrbl C0=Crbl
xgc_0_1 wwl_0_1 wbl_0_1 rwl_0_1 rbl_0_1 sn_0_1 wos_ros_gc
xrc_wwl_0_1 wwl_0_0 wwl_0_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_1 wbl_1 wbl_0_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_1 rwl_0_0 rwl_0_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_1 rbl_1 rbl_0_1 rc_unit R0=Rrbl C0=Crbl
xgc_0_2 wwl_0_2 wbl_0_2 rwl_0_2 rbl_0_2 sn_0_2 wos_ros_gc
xrc_wwl_0_2 wwl_0_1 wwl_0_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_2 wbl_2 wbl_0_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_2 rwl_0_1 rwl_0_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_2 rbl_2 rbl_0_2 rc_unit R0=Rrbl C0=Crbl
xgc_0_3 wwl_0_3 wbl_0_3 rwl_0_3 rbl_0_3 sn_0_3 wos_ros_gc
xrc_wwl_0_3 wwl_0_2 wwl_0_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_3 wbl_3 wbl_0_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_3 rwl_0_2 rwl_0_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_3 rbl_3 rbl_0_3 rc_unit R0=Rrbl C0=Crbl
xgc_0_4 wwl_0_4 wbl_0_4 rwl_0_4 rbl_0_4 sn_0_4 wos_ros_gc
xrc_wwl_0_4 wwl_0_3 wwl_0_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_4 wbl_4 wbl_0_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_4 rwl_0_3 rwl_0_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_4 rbl_4 rbl_0_4 rc_unit R0=Rrbl C0=Crbl
xgc_0_5 wwl_0_5 wbl_0_5 rwl_0_5 rbl_0_5 sn_0_5 wos_ros_gc
xrc_wwl_0_5 wwl_0_4 wwl_0_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_5 wbl_5 wbl_0_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_5 rwl_0_4 rwl_0_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_5 rbl_5 rbl_0_5 rc_unit R0=Rrbl C0=Crbl
xgc_0_6 wwl_0_6 wbl_0_6 rwl_0_6 rbl_0_6 sn_0_6 wos_ros_gc
xrc_wwl_0_6 wwl_0_5 wwl_0_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_6 wbl_6 wbl_0_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_6 rwl_0_5 rwl_0_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_6 rbl_6 rbl_0_6 rc_unit R0=Rrbl C0=Crbl
xgc_0_7 wwl_0_7 wbl_0_7 rwl_0_7 rbl_0_7 sn_0_7 wos_ros_gc
xrc_wwl_0_7 wwl_0_6 wwl_0_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_7 wbl_7 wbl_0_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_7 rwl_0_6 rwl_0_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_7 rbl_7 rbl_0_7 rc_unit R0=Rrbl C0=Crbl
xgc_0_8 wwl_0_8 wbl_0_8 rwl_0_8 rbl_0_8 sn_0_8 wos_ros_gc
xrc_wwl_0_8 wwl_0_7 wwl_0_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_8 wbl_8 wbl_0_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_8 rwl_0_7 rwl_0_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_8 rbl_8 rbl_0_8 rc_unit R0=Rrbl C0=Crbl
xgc_0_9 wwl_0_9 wbl_0_9 rwl_0_9 rbl_0_9 sn_0_9 wos_ros_gc
xrc_wwl_0_9 wwl_0_8 wwl_0_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_9 wbl_9 wbl_0_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_9 rwl_0_8 rwl_0_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_9 rbl_9 rbl_0_9 rc_unit R0=Rrbl C0=Crbl
xgc_0_10 wwl_0_10 wbl_0_10 rwl_0_10 rbl_0_10 sn_0_10 wos_ros_gc
xrc_wwl_0_10 wwl_0_9 wwl_0_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_10 wbl_10 wbl_0_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_10 rwl_0_9 rwl_0_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_10 rbl_10 rbl_0_10 rc_unit R0=Rrbl C0=Crbl
xgc_0_11 wwl_0_11 wbl_0_11 rwl_0_11 rbl_0_11 sn_0_11 wos_ros_gc
xrc_wwl_0_11 wwl_0_10 wwl_0_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_11 wbl_11 wbl_0_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_11 rwl_0_10 rwl_0_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_11 rbl_11 rbl_0_11 rc_unit R0=Rrbl C0=Crbl
xgc_0_12 wwl_0_12 wbl_0_12 rwl_0_12 rbl_0_12 sn_0_12 wos_ros_gc
xrc_wwl_0_12 wwl_0_11 wwl_0_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_12 wbl_12 wbl_0_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_12 rwl_0_11 rwl_0_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_12 rbl_12 rbl_0_12 rc_unit R0=Rrbl C0=Crbl
xgc_0_13 wwl_0_13 wbl_0_13 rwl_0_13 rbl_0_13 sn_0_13 wos_ros_gc
xrc_wwl_0_13 wwl_0_12 wwl_0_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_13 wbl_13 wbl_0_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_13 rwl_0_12 rwl_0_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_13 rbl_13 rbl_0_13 rc_unit R0=Rrbl C0=Crbl
xgc_0_14 wwl_0_14 wbl_0_14 rwl_0_14 rbl_0_14 sn_0_14 wos_ros_gc
xrc_wwl_0_14 wwl_0_13 wwl_0_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_14 wbl_14 wbl_0_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_14 rwl_0_13 rwl_0_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_14 rbl_14 rbl_0_14 rc_unit R0=Rrbl C0=Crbl
xgc_0_15 wwl_0_15 wbl_0_15 rwl_0_15 rbl_0_15 sn_0_15 wos_ros_gc
xrc_wwl_0_15 wwl_0_14 wwl_0_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_15 wbl_15 wbl_0_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_15 rwl_0_14 rwl_0_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_15 rbl_15 rbl_0_15 rc_unit R0=Rrbl C0=Crbl
xgc_0_16 wwl_0_16 wbl_0_16 rwl_0_16 rbl_0_16 sn_0_16 wos_ros_gc
xrc_wwl_0_16 wwl_0_15 wwl_0_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_16 wbl_16 wbl_0_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_16 rwl_0_15 rwl_0_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_16 rbl_16 rbl_0_16 rc_unit R0=Rrbl C0=Crbl
xgc_0_17 wwl_0_17 wbl_0_17 rwl_0_17 rbl_0_17 sn_0_17 wos_ros_gc
xrc_wwl_0_17 wwl_0_16 wwl_0_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_17 wbl_17 wbl_0_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_17 rwl_0_16 rwl_0_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_17 rbl_17 rbl_0_17 rc_unit R0=Rrbl C0=Crbl
xgc_0_18 wwl_0_18 wbl_0_18 rwl_0_18 rbl_0_18 sn_0_18 wos_ros_gc
xrc_wwl_0_18 wwl_0_17 wwl_0_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_18 wbl_18 wbl_0_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_18 rwl_0_17 rwl_0_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_18 rbl_18 rbl_0_18 rc_unit R0=Rrbl C0=Crbl
xgc_0_19 wwl_0_19 wbl_0_19 rwl_0_19 rbl_0_19 sn_0_19 wos_ros_gc
xrc_wwl_0_19 wwl_0_18 wwl_0_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_19 wbl_19 wbl_0_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_19 rwl_0_18 rwl_0_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_19 rbl_19 rbl_0_19 rc_unit R0=Rrbl C0=Crbl
xgc_0_20 wwl_0_20 wbl_0_20 rwl_0_20 rbl_0_20 sn_0_20 wos_ros_gc
xrc_wwl_0_20 wwl_0_19 wwl_0_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_20 wbl_20 wbl_0_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_20 rwl_0_19 rwl_0_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_20 rbl_20 rbl_0_20 rc_unit R0=Rrbl C0=Crbl
xgc_0_21 wwl_0_21 wbl_0_21 rwl_0_21 rbl_0_21 sn_0_21 wos_ros_gc
xrc_wwl_0_21 wwl_0_20 wwl_0_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_21 wbl_21 wbl_0_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_21 rwl_0_20 rwl_0_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_21 rbl_21 rbl_0_21 rc_unit R0=Rrbl C0=Crbl
xgc_0_22 wwl_0_22 wbl_0_22 rwl_0_22 rbl_0_22 sn_0_22 wos_ros_gc
xrc_wwl_0_22 wwl_0_21 wwl_0_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_22 wbl_22 wbl_0_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_22 rwl_0_21 rwl_0_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_22 rbl_22 rbl_0_22 rc_unit R0=Rrbl C0=Crbl
xgc_0_23 wwl_0_23 wbl_0_23 rwl_0_23 rbl_0_23 sn_0_23 wos_ros_gc
xrc_wwl_0_23 wwl_0_22 wwl_0_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_23 wbl_23 wbl_0_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_23 rwl_0_22 rwl_0_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_23 rbl_23 rbl_0_23 rc_unit R0=Rrbl C0=Crbl
xgc_0_24 wwl_0_24 wbl_0_24 rwl_0_24 rbl_0_24 sn_0_24 wos_ros_gc
xrc_wwl_0_24 wwl_0_23 wwl_0_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_24 wbl_24 wbl_0_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_24 rwl_0_23 rwl_0_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_24 rbl_24 rbl_0_24 rc_unit R0=Rrbl C0=Crbl
xgc_0_25 wwl_0_25 wbl_0_25 rwl_0_25 rbl_0_25 sn_0_25 wos_ros_gc
xrc_wwl_0_25 wwl_0_24 wwl_0_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_25 wbl_25 wbl_0_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_25 rwl_0_24 rwl_0_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_25 rbl_25 rbl_0_25 rc_unit R0=Rrbl C0=Crbl
xgc_0_26 wwl_0_26 wbl_0_26 rwl_0_26 rbl_0_26 sn_0_26 wos_ros_gc
xrc_wwl_0_26 wwl_0_25 wwl_0_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_26 wbl_26 wbl_0_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_26 rwl_0_25 rwl_0_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_26 rbl_26 rbl_0_26 rc_unit R0=Rrbl C0=Crbl
xgc_0_27 wwl_0_27 wbl_0_27 rwl_0_27 rbl_0_27 sn_0_27 wos_ros_gc
xrc_wwl_0_27 wwl_0_26 wwl_0_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_27 wbl_27 wbl_0_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_27 rwl_0_26 rwl_0_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_27 rbl_27 rbl_0_27 rc_unit R0=Rrbl C0=Crbl
xgc_0_28 wwl_0_28 wbl_0_28 rwl_0_28 rbl_0_28 sn_0_28 wos_ros_gc
xrc_wwl_0_28 wwl_0_27 wwl_0_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_28 wbl_28 wbl_0_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_28 rwl_0_27 rwl_0_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_28 rbl_28 rbl_0_28 rc_unit R0=Rrbl C0=Crbl
xgc_0_29 wwl_0_29 wbl_0_29 rwl_0_29 rbl_0_29 sn_0_29 wos_ros_gc
xrc_wwl_0_29 wwl_0_28 wwl_0_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_29 wbl_29 wbl_0_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_29 rwl_0_28 rwl_0_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_29 rbl_29 rbl_0_29 rc_unit R0=Rrbl C0=Crbl
xgc_0_30 wwl_0_30 wbl_0_30 rwl_0_30 rbl_0_30 sn_0_30 wos_ros_gc
xrc_wwl_0_30 wwl_0_29 wwl_0_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_30 wbl_30 wbl_0_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_30 rwl_0_29 rwl_0_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_30 rbl_30 rbl_0_30 rc_unit R0=Rrbl C0=Crbl
xgc_0_31 wwl_0_31 wbl_0_31 rwl_0_31 rbl_0_31 sn_0_31 wos_ros_gc
xrc_wwl_0_31 wwl_0_30 wwl_0_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_0_31 wbl_31 wbl_0_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_0_31 rwl_0_30 rwl_0_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_0_31 rbl_31 rbl_0_31 rc_unit R0=Rrbl C0=Crbl
xgc_1_0 wwl_1_0 wbl_1_0 rwl_1_0 rbl_1_0 sn_1_0 wos_ros_gc
xrc_wwl_1_0 wwl_1 wwl_1_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_0 wbl_0_0 wbl_1_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_0 rwl_1 rwl_1_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_0 rbl_0_0 rbl_1_0 rc_unit R0=Rrbl C0=Crbl
xgc_1_1 wwl_1_1 wbl_1_1 rwl_1_1 rbl_1_1 sn_1_1 wos_ros_gc
xrc_wwl_1_1 wwl_1_0 wwl_1_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_1 wbl_0_1 wbl_1_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_1 rwl_1_0 rwl_1_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_1 rbl_0_1 rbl_1_1 rc_unit R0=Rrbl C0=Crbl
xgc_1_2 wwl_1_2 wbl_1_2 rwl_1_2 rbl_1_2 sn_1_2 wos_ros_gc
xrc_wwl_1_2 wwl_1_1 wwl_1_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_2 wbl_0_2 wbl_1_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_2 rwl_1_1 rwl_1_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_2 rbl_0_2 rbl_1_2 rc_unit R0=Rrbl C0=Crbl
xgc_1_3 wwl_1_3 wbl_1_3 rwl_1_3 rbl_1_3 sn_1_3 wos_ros_gc
xrc_wwl_1_3 wwl_1_2 wwl_1_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_3 wbl_0_3 wbl_1_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_3 rwl_1_2 rwl_1_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_3 rbl_0_3 rbl_1_3 rc_unit R0=Rrbl C0=Crbl
xgc_1_4 wwl_1_4 wbl_1_4 rwl_1_4 rbl_1_4 sn_1_4 wos_ros_gc
xrc_wwl_1_4 wwl_1_3 wwl_1_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_4 wbl_0_4 wbl_1_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_4 rwl_1_3 rwl_1_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_4 rbl_0_4 rbl_1_4 rc_unit R0=Rrbl C0=Crbl
xgc_1_5 wwl_1_5 wbl_1_5 rwl_1_5 rbl_1_5 sn_1_5 wos_ros_gc
xrc_wwl_1_5 wwl_1_4 wwl_1_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_5 wbl_0_5 wbl_1_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_5 rwl_1_4 rwl_1_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_5 rbl_0_5 rbl_1_5 rc_unit R0=Rrbl C0=Crbl
xgc_1_6 wwl_1_6 wbl_1_6 rwl_1_6 rbl_1_6 sn_1_6 wos_ros_gc
xrc_wwl_1_6 wwl_1_5 wwl_1_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_6 wbl_0_6 wbl_1_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_6 rwl_1_5 rwl_1_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_6 rbl_0_6 rbl_1_6 rc_unit R0=Rrbl C0=Crbl
xgc_1_7 wwl_1_7 wbl_1_7 rwl_1_7 rbl_1_7 sn_1_7 wos_ros_gc
xrc_wwl_1_7 wwl_1_6 wwl_1_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_7 wbl_0_7 wbl_1_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_7 rwl_1_6 rwl_1_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_7 rbl_0_7 rbl_1_7 rc_unit R0=Rrbl C0=Crbl
xgc_1_8 wwl_1_8 wbl_1_8 rwl_1_8 rbl_1_8 sn_1_8 wos_ros_gc
xrc_wwl_1_8 wwl_1_7 wwl_1_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_8 wbl_0_8 wbl_1_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_8 rwl_1_7 rwl_1_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_8 rbl_0_8 rbl_1_8 rc_unit R0=Rrbl C0=Crbl
xgc_1_9 wwl_1_9 wbl_1_9 rwl_1_9 rbl_1_9 sn_1_9 wos_ros_gc
xrc_wwl_1_9 wwl_1_8 wwl_1_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_9 wbl_0_9 wbl_1_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_9 rwl_1_8 rwl_1_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_9 rbl_0_9 rbl_1_9 rc_unit R0=Rrbl C0=Crbl
xgc_1_10 wwl_1_10 wbl_1_10 rwl_1_10 rbl_1_10 sn_1_10 wos_ros_gc
xrc_wwl_1_10 wwl_1_9 wwl_1_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_10 wbl_0_10 wbl_1_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_10 rwl_1_9 rwl_1_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_10 rbl_0_10 rbl_1_10 rc_unit R0=Rrbl C0=Crbl
xgc_1_11 wwl_1_11 wbl_1_11 rwl_1_11 rbl_1_11 sn_1_11 wos_ros_gc
xrc_wwl_1_11 wwl_1_10 wwl_1_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_11 wbl_0_11 wbl_1_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_11 rwl_1_10 rwl_1_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_11 rbl_0_11 rbl_1_11 rc_unit R0=Rrbl C0=Crbl
xgc_1_12 wwl_1_12 wbl_1_12 rwl_1_12 rbl_1_12 sn_1_12 wos_ros_gc
xrc_wwl_1_12 wwl_1_11 wwl_1_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_12 wbl_0_12 wbl_1_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_12 rwl_1_11 rwl_1_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_12 rbl_0_12 rbl_1_12 rc_unit R0=Rrbl C0=Crbl
xgc_1_13 wwl_1_13 wbl_1_13 rwl_1_13 rbl_1_13 sn_1_13 wos_ros_gc
xrc_wwl_1_13 wwl_1_12 wwl_1_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_13 wbl_0_13 wbl_1_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_13 rwl_1_12 rwl_1_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_13 rbl_0_13 rbl_1_13 rc_unit R0=Rrbl C0=Crbl
xgc_1_14 wwl_1_14 wbl_1_14 rwl_1_14 rbl_1_14 sn_1_14 wos_ros_gc
xrc_wwl_1_14 wwl_1_13 wwl_1_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_14 wbl_0_14 wbl_1_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_14 rwl_1_13 rwl_1_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_14 rbl_0_14 rbl_1_14 rc_unit R0=Rrbl C0=Crbl
xgc_1_15 wwl_1_15 wbl_1_15 rwl_1_15 rbl_1_15 sn_1_15 wos_ros_gc
xrc_wwl_1_15 wwl_1_14 wwl_1_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_15 wbl_0_15 wbl_1_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_15 rwl_1_14 rwl_1_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_15 rbl_0_15 rbl_1_15 rc_unit R0=Rrbl C0=Crbl
xgc_1_16 wwl_1_16 wbl_1_16 rwl_1_16 rbl_1_16 sn_1_16 wos_ros_gc
xrc_wwl_1_16 wwl_1_15 wwl_1_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_16 wbl_0_16 wbl_1_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_16 rwl_1_15 rwl_1_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_16 rbl_0_16 rbl_1_16 rc_unit R0=Rrbl C0=Crbl
xgc_1_17 wwl_1_17 wbl_1_17 rwl_1_17 rbl_1_17 sn_1_17 wos_ros_gc
xrc_wwl_1_17 wwl_1_16 wwl_1_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_17 wbl_0_17 wbl_1_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_17 rwl_1_16 rwl_1_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_17 rbl_0_17 rbl_1_17 rc_unit R0=Rrbl C0=Crbl
xgc_1_18 wwl_1_18 wbl_1_18 rwl_1_18 rbl_1_18 sn_1_18 wos_ros_gc
xrc_wwl_1_18 wwl_1_17 wwl_1_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_18 wbl_0_18 wbl_1_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_18 rwl_1_17 rwl_1_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_18 rbl_0_18 rbl_1_18 rc_unit R0=Rrbl C0=Crbl
xgc_1_19 wwl_1_19 wbl_1_19 rwl_1_19 rbl_1_19 sn_1_19 wos_ros_gc
xrc_wwl_1_19 wwl_1_18 wwl_1_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_19 wbl_0_19 wbl_1_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_19 rwl_1_18 rwl_1_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_19 rbl_0_19 rbl_1_19 rc_unit R0=Rrbl C0=Crbl
xgc_1_20 wwl_1_20 wbl_1_20 rwl_1_20 rbl_1_20 sn_1_20 wos_ros_gc
xrc_wwl_1_20 wwl_1_19 wwl_1_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_20 wbl_0_20 wbl_1_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_20 rwl_1_19 rwl_1_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_20 rbl_0_20 rbl_1_20 rc_unit R0=Rrbl C0=Crbl
xgc_1_21 wwl_1_21 wbl_1_21 rwl_1_21 rbl_1_21 sn_1_21 wos_ros_gc
xrc_wwl_1_21 wwl_1_20 wwl_1_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_21 wbl_0_21 wbl_1_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_21 rwl_1_20 rwl_1_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_21 rbl_0_21 rbl_1_21 rc_unit R0=Rrbl C0=Crbl
xgc_1_22 wwl_1_22 wbl_1_22 rwl_1_22 rbl_1_22 sn_1_22 wos_ros_gc
xrc_wwl_1_22 wwl_1_21 wwl_1_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_22 wbl_0_22 wbl_1_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_22 rwl_1_21 rwl_1_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_22 rbl_0_22 rbl_1_22 rc_unit R0=Rrbl C0=Crbl
xgc_1_23 wwl_1_23 wbl_1_23 rwl_1_23 rbl_1_23 sn_1_23 wos_ros_gc
xrc_wwl_1_23 wwl_1_22 wwl_1_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_23 wbl_0_23 wbl_1_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_23 rwl_1_22 rwl_1_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_23 rbl_0_23 rbl_1_23 rc_unit R0=Rrbl C0=Crbl
xgc_1_24 wwl_1_24 wbl_1_24 rwl_1_24 rbl_1_24 sn_1_24 wos_ros_gc
xrc_wwl_1_24 wwl_1_23 wwl_1_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_24 wbl_0_24 wbl_1_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_24 rwl_1_23 rwl_1_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_24 rbl_0_24 rbl_1_24 rc_unit R0=Rrbl C0=Crbl
xgc_1_25 wwl_1_25 wbl_1_25 rwl_1_25 rbl_1_25 sn_1_25 wos_ros_gc
xrc_wwl_1_25 wwl_1_24 wwl_1_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_25 wbl_0_25 wbl_1_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_25 rwl_1_24 rwl_1_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_25 rbl_0_25 rbl_1_25 rc_unit R0=Rrbl C0=Crbl
xgc_1_26 wwl_1_26 wbl_1_26 rwl_1_26 rbl_1_26 sn_1_26 wos_ros_gc
xrc_wwl_1_26 wwl_1_25 wwl_1_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_26 wbl_0_26 wbl_1_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_26 rwl_1_25 rwl_1_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_26 rbl_0_26 rbl_1_26 rc_unit R0=Rrbl C0=Crbl
xgc_1_27 wwl_1_27 wbl_1_27 rwl_1_27 rbl_1_27 sn_1_27 wos_ros_gc
xrc_wwl_1_27 wwl_1_26 wwl_1_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_27 wbl_0_27 wbl_1_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_27 rwl_1_26 rwl_1_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_27 rbl_0_27 rbl_1_27 rc_unit R0=Rrbl C0=Crbl
xgc_1_28 wwl_1_28 wbl_1_28 rwl_1_28 rbl_1_28 sn_1_28 wos_ros_gc
xrc_wwl_1_28 wwl_1_27 wwl_1_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_28 wbl_0_28 wbl_1_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_28 rwl_1_27 rwl_1_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_28 rbl_0_28 rbl_1_28 rc_unit R0=Rrbl C0=Crbl
xgc_1_29 wwl_1_29 wbl_1_29 rwl_1_29 rbl_1_29 sn_1_29 wos_ros_gc
xrc_wwl_1_29 wwl_1_28 wwl_1_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_29 wbl_0_29 wbl_1_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_29 rwl_1_28 rwl_1_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_29 rbl_0_29 rbl_1_29 rc_unit R0=Rrbl C0=Crbl
xgc_1_30 wwl_1_30 wbl_1_30 rwl_1_30 rbl_1_30 sn_1_30 wos_ros_gc
xrc_wwl_1_30 wwl_1_29 wwl_1_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_30 wbl_0_30 wbl_1_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_30 rwl_1_29 rwl_1_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_30 rbl_0_30 rbl_1_30 rc_unit R0=Rrbl C0=Crbl
xgc_1_31 wwl_1_31 wbl_1_31 rwl_1_31 rbl_1_31 sn_1_31 wos_ros_gc
xrc_wwl_1_31 wwl_1_30 wwl_1_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_1_31 wbl_0_31 wbl_1_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_1_31 rwl_1_30 rwl_1_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_1_31 rbl_0_31 rbl_1_31 rc_unit R0=Rrbl C0=Crbl
xgc_2_0 wwl_2_0 wbl_2_0 rwl_2_0 rbl_2_0 sn_2_0 wos_ros_gc
xrc_wwl_2_0 wwl_2 wwl_2_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_0 wbl_1_0 wbl_2_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_0 rwl_2 rwl_2_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_0 rbl_1_0 rbl_2_0 rc_unit R0=Rrbl C0=Crbl
xgc_2_1 wwl_2_1 wbl_2_1 rwl_2_1 rbl_2_1 sn_2_1 wos_ros_gc
xrc_wwl_2_1 wwl_2_0 wwl_2_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_1 wbl_1_1 wbl_2_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_1 rwl_2_0 rwl_2_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_1 rbl_1_1 rbl_2_1 rc_unit R0=Rrbl C0=Crbl
xgc_2_2 wwl_2_2 wbl_2_2 rwl_2_2 rbl_2_2 sn_2_2 wos_ros_gc
xrc_wwl_2_2 wwl_2_1 wwl_2_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_2 wbl_1_2 wbl_2_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_2 rwl_2_1 rwl_2_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_2 rbl_1_2 rbl_2_2 rc_unit R0=Rrbl C0=Crbl
xgc_2_3 wwl_2_3 wbl_2_3 rwl_2_3 rbl_2_3 sn_2_3 wos_ros_gc
xrc_wwl_2_3 wwl_2_2 wwl_2_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_3 wbl_1_3 wbl_2_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_3 rwl_2_2 rwl_2_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_3 rbl_1_3 rbl_2_3 rc_unit R0=Rrbl C0=Crbl
xgc_2_4 wwl_2_4 wbl_2_4 rwl_2_4 rbl_2_4 sn_2_4 wos_ros_gc
xrc_wwl_2_4 wwl_2_3 wwl_2_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_4 wbl_1_4 wbl_2_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_4 rwl_2_3 rwl_2_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_4 rbl_1_4 rbl_2_4 rc_unit R0=Rrbl C0=Crbl
xgc_2_5 wwl_2_5 wbl_2_5 rwl_2_5 rbl_2_5 sn_2_5 wos_ros_gc
xrc_wwl_2_5 wwl_2_4 wwl_2_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_5 wbl_1_5 wbl_2_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_5 rwl_2_4 rwl_2_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_5 rbl_1_5 rbl_2_5 rc_unit R0=Rrbl C0=Crbl
xgc_2_6 wwl_2_6 wbl_2_6 rwl_2_6 rbl_2_6 sn_2_6 wos_ros_gc
xrc_wwl_2_6 wwl_2_5 wwl_2_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_6 wbl_1_6 wbl_2_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_6 rwl_2_5 rwl_2_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_6 rbl_1_6 rbl_2_6 rc_unit R0=Rrbl C0=Crbl
xgc_2_7 wwl_2_7 wbl_2_7 rwl_2_7 rbl_2_7 sn_2_7 wos_ros_gc
xrc_wwl_2_7 wwl_2_6 wwl_2_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_7 wbl_1_7 wbl_2_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_7 rwl_2_6 rwl_2_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_7 rbl_1_7 rbl_2_7 rc_unit R0=Rrbl C0=Crbl
xgc_2_8 wwl_2_8 wbl_2_8 rwl_2_8 rbl_2_8 sn_2_8 wos_ros_gc
xrc_wwl_2_8 wwl_2_7 wwl_2_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_8 wbl_1_8 wbl_2_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_8 rwl_2_7 rwl_2_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_8 rbl_1_8 rbl_2_8 rc_unit R0=Rrbl C0=Crbl
xgc_2_9 wwl_2_9 wbl_2_9 rwl_2_9 rbl_2_9 sn_2_9 wos_ros_gc
xrc_wwl_2_9 wwl_2_8 wwl_2_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_9 wbl_1_9 wbl_2_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_9 rwl_2_8 rwl_2_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_9 rbl_1_9 rbl_2_9 rc_unit R0=Rrbl C0=Crbl
xgc_2_10 wwl_2_10 wbl_2_10 rwl_2_10 rbl_2_10 sn_2_10 wos_ros_gc
xrc_wwl_2_10 wwl_2_9 wwl_2_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_10 wbl_1_10 wbl_2_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_10 rwl_2_9 rwl_2_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_10 rbl_1_10 rbl_2_10 rc_unit R0=Rrbl C0=Crbl
xgc_2_11 wwl_2_11 wbl_2_11 rwl_2_11 rbl_2_11 sn_2_11 wos_ros_gc
xrc_wwl_2_11 wwl_2_10 wwl_2_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_11 wbl_1_11 wbl_2_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_11 rwl_2_10 rwl_2_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_11 rbl_1_11 rbl_2_11 rc_unit R0=Rrbl C0=Crbl
xgc_2_12 wwl_2_12 wbl_2_12 rwl_2_12 rbl_2_12 sn_2_12 wos_ros_gc
xrc_wwl_2_12 wwl_2_11 wwl_2_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_12 wbl_1_12 wbl_2_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_12 rwl_2_11 rwl_2_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_12 rbl_1_12 rbl_2_12 rc_unit R0=Rrbl C0=Crbl
xgc_2_13 wwl_2_13 wbl_2_13 rwl_2_13 rbl_2_13 sn_2_13 wos_ros_gc
xrc_wwl_2_13 wwl_2_12 wwl_2_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_13 wbl_1_13 wbl_2_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_13 rwl_2_12 rwl_2_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_13 rbl_1_13 rbl_2_13 rc_unit R0=Rrbl C0=Crbl
xgc_2_14 wwl_2_14 wbl_2_14 rwl_2_14 rbl_2_14 sn_2_14 wos_ros_gc
xrc_wwl_2_14 wwl_2_13 wwl_2_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_14 wbl_1_14 wbl_2_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_14 rwl_2_13 rwl_2_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_14 rbl_1_14 rbl_2_14 rc_unit R0=Rrbl C0=Crbl
xgc_2_15 wwl_2_15 wbl_2_15 rwl_2_15 rbl_2_15 sn_2_15 wos_ros_gc
xrc_wwl_2_15 wwl_2_14 wwl_2_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_15 wbl_1_15 wbl_2_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_15 rwl_2_14 rwl_2_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_15 rbl_1_15 rbl_2_15 rc_unit R0=Rrbl C0=Crbl
xgc_2_16 wwl_2_16 wbl_2_16 rwl_2_16 rbl_2_16 sn_2_16 wos_ros_gc
xrc_wwl_2_16 wwl_2_15 wwl_2_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_16 wbl_1_16 wbl_2_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_16 rwl_2_15 rwl_2_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_16 rbl_1_16 rbl_2_16 rc_unit R0=Rrbl C0=Crbl
xgc_2_17 wwl_2_17 wbl_2_17 rwl_2_17 rbl_2_17 sn_2_17 wos_ros_gc
xrc_wwl_2_17 wwl_2_16 wwl_2_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_17 wbl_1_17 wbl_2_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_17 rwl_2_16 rwl_2_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_17 rbl_1_17 rbl_2_17 rc_unit R0=Rrbl C0=Crbl
xgc_2_18 wwl_2_18 wbl_2_18 rwl_2_18 rbl_2_18 sn_2_18 wos_ros_gc
xrc_wwl_2_18 wwl_2_17 wwl_2_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_18 wbl_1_18 wbl_2_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_18 rwl_2_17 rwl_2_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_18 rbl_1_18 rbl_2_18 rc_unit R0=Rrbl C0=Crbl
xgc_2_19 wwl_2_19 wbl_2_19 rwl_2_19 rbl_2_19 sn_2_19 wos_ros_gc
xrc_wwl_2_19 wwl_2_18 wwl_2_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_19 wbl_1_19 wbl_2_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_19 rwl_2_18 rwl_2_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_19 rbl_1_19 rbl_2_19 rc_unit R0=Rrbl C0=Crbl
xgc_2_20 wwl_2_20 wbl_2_20 rwl_2_20 rbl_2_20 sn_2_20 wos_ros_gc
xrc_wwl_2_20 wwl_2_19 wwl_2_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_20 wbl_1_20 wbl_2_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_20 rwl_2_19 rwl_2_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_20 rbl_1_20 rbl_2_20 rc_unit R0=Rrbl C0=Crbl
xgc_2_21 wwl_2_21 wbl_2_21 rwl_2_21 rbl_2_21 sn_2_21 wos_ros_gc
xrc_wwl_2_21 wwl_2_20 wwl_2_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_21 wbl_1_21 wbl_2_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_21 rwl_2_20 rwl_2_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_21 rbl_1_21 rbl_2_21 rc_unit R0=Rrbl C0=Crbl
xgc_2_22 wwl_2_22 wbl_2_22 rwl_2_22 rbl_2_22 sn_2_22 wos_ros_gc
xrc_wwl_2_22 wwl_2_21 wwl_2_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_22 wbl_1_22 wbl_2_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_22 rwl_2_21 rwl_2_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_22 rbl_1_22 rbl_2_22 rc_unit R0=Rrbl C0=Crbl
xgc_2_23 wwl_2_23 wbl_2_23 rwl_2_23 rbl_2_23 sn_2_23 wos_ros_gc
xrc_wwl_2_23 wwl_2_22 wwl_2_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_23 wbl_1_23 wbl_2_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_23 rwl_2_22 rwl_2_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_23 rbl_1_23 rbl_2_23 rc_unit R0=Rrbl C0=Crbl
xgc_2_24 wwl_2_24 wbl_2_24 rwl_2_24 rbl_2_24 sn_2_24 wos_ros_gc
xrc_wwl_2_24 wwl_2_23 wwl_2_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_24 wbl_1_24 wbl_2_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_24 rwl_2_23 rwl_2_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_24 rbl_1_24 rbl_2_24 rc_unit R0=Rrbl C0=Crbl
xgc_2_25 wwl_2_25 wbl_2_25 rwl_2_25 rbl_2_25 sn_2_25 wos_ros_gc
xrc_wwl_2_25 wwl_2_24 wwl_2_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_25 wbl_1_25 wbl_2_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_25 rwl_2_24 rwl_2_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_25 rbl_1_25 rbl_2_25 rc_unit R0=Rrbl C0=Crbl
xgc_2_26 wwl_2_26 wbl_2_26 rwl_2_26 rbl_2_26 sn_2_26 wos_ros_gc
xrc_wwl_2_26 wwl_2_25 wwl_2_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_26 wbl_1_26 wbl_2_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_26 rwl_2_25 rwl_2_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_26 rbl_1_26 rbl_2_26 rc_unit R0=Rrbl C0=Crbl
xgc_2_27 wwl_2_27 wbl_2_27 rwl_2_27 rbl_2_27 sn_2_27 wos_ros_gc
xrc_wwl_2_27 wwl_2_26 wwl_2_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_27 wbl_1_27 wbl_2_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_27 rwl_2_26 rwl_2_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_27 rbl_1_27 rbl_2_27 rc_unit R0=Rrbl C0=Crbl
xgc_2_28 wwl_2_28 wbl_2_28 rwl_2_28 rbl_2_28 sn_2_28 wos_ros_gc
xrc_wwl_2_28 wwl_2_27 wwl_2_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_28 wbl_1_28 wbl_2_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_28 rwl_2_27 rwl_2_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_28 rbl_1_28 rbl_2_28 rc_unit R0=Rrbl C0=Crbl
xgc_2_29 wwl_2_29 wbl_2_29 rwl_2_29 rbl_2_29 sn_2_29 wos_ros_gc
xrc_wwl_2_29 wwl_2_28 wwl_2_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_29 wbl_1_29 wbl_2_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_29 rwl_2_28 rwl_2_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_29 rbl_1_29 rbl_2_29 rc_unit R0=Rrbl C0=Crbl
xgc_2_30 wwl_2_30 wbl_2_30 rwl_2_30 rbl_2_30 sn_2_30 wos_ros_gc
xrc_wwl_2_30 wwl_2_29 wwl_2_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_30 wbl_1_30 wbl_2_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_30 rwl_2_29 rwl_2_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_30 rbl_1_30 rbl_2_30 rc_unit R0=Rrbl C0=Crbl
xgc_2_31 wwl_2_31 wbl_2_31 rwl_2_31 rbl_2_31 sn_2_31 wos_ros_gc
xrc_wwl_2_31 wwl_2_30 wwl_2_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_2_31 wbl_1_31 wbl_2_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_2_31 rwl_2_30 rwl_2_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_2_31 rbl_1_31 rbl_2_31 rc_unit R0=Rrbl C0=Crbl
xgc_3_0 wwl_3_0 wbl_3_0 rwl_3_0 rbl_3_0 sn_3_0 wos_ros_gc
xrc_wwl_3_0 wwl_3 wwl_3_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_0 wbl_2_0 wbl_3_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_0 rwl_3 rwl_3_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_0 rbl_2_0 rbl_3_0 rc_unit R0=Rrbl C0=Crbl
xgc_3_1 wwl_3_1 wbl_3_1 rwl_3_1 rbl_3_1 sn_3_1 wos_ros_gc
xrc_wwl_3_1 wwl_3_0 wwl_3_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_1 wbl_2_1 wbl_3_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_1 rwl_3_0 rwl_3_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_1 rbl_2_1 rbl_3_1 rc_unit R0=Rrbl C0=Crbl
xgc_3_2 wwl_3_2 wbl_3_2 rwl_3_2 rbl_3_2 sn_3_2 wos_ros_gc
xrc_wwl_3_2 wwl_3_1 wwl_3_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_2 wbl_2_2 wbl_3_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_2 rwl_3_1 rwl_3_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_2 rbl_2_2 rbl_3_2 rc_unit R0=Rrbl C0=Crbl
xgc_3_3 wwl_3_3 wbl_3_3 rwl_3_3 rbl_3_3 sn_3_3 wos_ros_gc
xrc_wwl_3_3 wwl_3_2 wwl_3_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_3 wbl_2_3 wbl_3_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_3 rwl_3_2 rwl_3_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_3 rbl_2_3 rbl_3_3 rc_unit R0=Rrbl C0=Crbl
xgc_3_4 wwl_3_4 wbl_3_4 rwl_3_4 rbl_3_4 sn_3_4 wos_ros_gc
xrc_wwl_3_4 wwl_3_3 wwl_3_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_4 wbl_2_4 wbl_3_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_4 rwl_3_3 rwl_3_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_4 rbl_2_4 rbl_3_4 rc_unit R0=Rrbl C0=Crbl
xgc_3_5 wwl_3_5 wbl_3_5 rwl_3_5 rbl_3_5 sn_3_5 wos_ros_gc
xrc_wwl_3_5 wwl_3_4 wwl_3_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_5 wbl_2_5 wbl_3_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_5 rwl_3_4 rwl_3_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_5 rbl_2_5 rbl_3_5 rc_unit R0=Rrbl C0=Crbl
xgc_3_6 wwl_3_6 wbl_3_6 rwl_3_6 rbl_3_6 sn_3_6 wos_ros_gc
xrc_wwl_3_6 wwl_3_5 wwl_3_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_6 wbl_2_6 wbl_3_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_6 rwl_3_5 rwl_3_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_6 rbl_2_6 rbl_3_6 rc_unit R0=Rrbl C0=Crbl
xgc_3_7 wwl_3_7 wbl_3_7 rwl_3_7 rbl_3_7 sn_3_7 wos_ros_gc
xrc_wwl_3_7 wwl_3_6 wwl_3_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_7 wbl_2_7 wbl_3_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_7 rwl_3_6 rwl_3_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_7 rbl_2_7 rbl_3_7 rc_unit R0=Rrbl C0=Crbl
xgc_3_8 wwl_3_8 wbl_3_8 rwl_3_8 rbl_3_8 sn_3_8 wos_ros_gc
xrc_wwl_3_8 wwl_3_7 wwl_3_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_8 wbl_2_8 wbl_3_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_8 rwl_3_7 rwl_3_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_8 rbl_2_8 rbl_3_8 rc_unit R0=Rrbl C0=Crbl
xgc_3_9 wwl_3_9 wbl_3_9 rwl_3_9 rbl_3_9 sn_3_9 wos_ros_gc
xrc_wwl_3_9 wwl_3_8 wwl_3_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_9 wbl_2_9 wbl_3_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_9 rwl_3_8 rwl_3_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_9 rbl_2_9 rbl_3_9 rc_unit R0=Rrbl C0=Crbl
xgc_3_10 wwl_3_10 wbl_3_10 rwl_3_10 rbl_3_10 sn_3_10 wos_ros_gc
xrc_wwl_3_10 wwl_3_9 wwl_3_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_10 wbl_2_10 wbl_3_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_10 rwl_3_9 rwl_3_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_10 rbl_2_10 rbl_3_10 rc_unit R0=Rrbl C0=Crbl
xgc_3_11 wwl_3_11 wbl_3_11 rwl_3_11 rbl_3_11 sn_3_11 wos_ros_gc
xrc_wwl_3_11 wwl_3_10 wwl_3_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_11 wbl_2_11 wbl_3_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_11 rwl_3_10 rwl_3_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_11 rbl_2_11 rbl_3_11 rc_unit R0=Rrbl C0=Crbl
xgc_3_12 wwl_3_12 wbl_3_12 rwl_3_12 rbl_3_12 sn_3_12 wos_ros_gc
xrc_wwl_3_12 wwl_3_11 wwl_3_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_12 wbl_2_12 wbl_3_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_12 rwl_3_11 rwl_3_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_12 rbl_2_12 rbl_3_12 rc_unit R0=Rrbl C0=Crbl
xgc_3_13 wwl_3_13 wbl_3_13 rwl_3_13 rbl_3_13 sn_3_13 wos_ros_gc
xrc_wwl_3_13 wwl_3_12 wwl_3_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_13 wbl_2_13 wbl_3_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_13 rwl_3_12 rwl_3_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_13 rbl_2_13 rbl_3_13 rc_unit R0=Rrbl C0=Crbl
xgc_3_14 wwl_3_14 wbl_3_14 rwl_3_14 rbl_3_14 sn_3_14 wos_ros_gc
xrc_wwl_3_14 wwl_3_13 wwl_3_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_14 wbl_2_14 wbl_3_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_14 rwl_3_13 rwl_3_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_14 rbl_2_14 rbl_3_14 rc_unit R0=Rrbl C0=Crbl
xgc_3_15 wwl_3_15 wbl_3_15 rwl_3_15 rbl_3_15 sn_3_15 wos_ros_gc
xrc_wwl_3_15 wwl_3_14 wwl_3_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_15 wbl_2_15 wbl_3_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_15 rwl_3_14 rwl_3_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_15 rbl_2_15 rbl_3_15 rc_unit R0=Rrbl C0=Crbl
xgc_3_16 wwl_3_16 wbl_3_16 rwl_3_16 rbl_3_16 sn_3_16 wos_ros_gc
xrc_wwl_3_16 wwl_3_15 wwl_3_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_16 wbl_2_16 wbl_3_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_16 rwl_3_15 rwl_3_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_16 rbl_2_16 rbl_3_16 rc_unit R0=Rrbl C0=Crbl
xgc_3_17 wwl_3_17 wbl_3_17 rwl_3_17 rbl_3_17 sn_3_17 wos_ros_gc
xrc_wwl_3_17 wwl_3_16 wwl_3_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_17 wbl_2_17 wbl_3_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_17 rwl_3_16 rwl_3_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_17 rbl_2_17 rbl_3_17 rc_unit R0=Rrbl C0=Crbl
xgc_3_18 wwl_3_18 wbl_3_18 rwl_3_18 rbl_3_18 sn_3_18 wos_ros_gc
xrc_wwl_3_18 wwl_3_17 wwl_3_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_18 wbl_2_18 wbl_3_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_18 rwl_3_17 rwl_3_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_18 rbl_2_18 rbl_3_18 rc_unit R0=Rrbl C0=Crbl
xgc_3_19 wwl_3_19 wbl_3_19 rwl_3_19 rbl_3_19 sn_3_19 wos_ros_gc
xrc_wwl_3_19 wwl_3_18 wwl_3_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_19 wbl_2_19 wbl_3_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_19 rwl_3_18 rwl_3_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_19 rbl_2_19 rbl_3_19 rc_unit R0=Rrbl C0=Crbl
xgc_3_20 wwl_3_20 wbl_3_20 rwl_3_20 rbl_3_20 sn_3_20 wos_ros_gc
xrc_wwl_3_20 wwl_3_19 wwl_3_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_20 wbl_2_20 wbl_3_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_20 rwl_3_19 rwl_3_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_20 rbl_2_20 rbl_3_20 rc_unit R0=Rrbl C0=Crbl
xgc_3_21 wwl_3_21 wbl_3_21 rwl_3_21 rbl_3_21 sn_3_21 wos_ros_gc
xrc_wwl_3_21 wwl_3_20 wwl_3_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_21 wbl_2_21 wbl_3_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_21 rwl_3_20 rwl_3_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_21 rbl_2_21 rbl_3_21 rc_unit R0=Rrbl C0=Crbl
xgc_3_22 wwl_3_22 wbl_3_22 rwl_3_22 rbl_3_22 sn_3_22 wos_ros_gc
xrc_wwl_3_22 wwl_3_21 wwl_3_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_22 wbl_2_22 wbl_3_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_22 rwl_3_21 rwl_3_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_22 rbl_2_22 rbl_3_22 rc_unit R0=Rrbl C0=Crbl
xgc_3_23 wwl_3_23 wbl_3_23 rwl_3_23 rbl_3_23 sn_3_23 wos_ros_gc
xrc_wwl_3_23 wwl_3_22 wwl_3_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_23 wbl_2_23 wbl_3_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_23 rwl_3_22 rwl_3_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_23 rbl_2_23 rbl_3_23 rc_unit R0=Rrbl C0=Crbl
xgc_3_24 wwl_3_24 wbl_3_24 rwl_3_24 rbl_3_24 sn_3_24 wos_ros_gc
xrc_wwl_3_24 wwl_3_23 wwl_3_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_24 wbl_2_24 wbl_3_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_24 rwl_3_23 rwl_3_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_24 rbl_2_24 rbl_3_24 rc_unit R0=Rrbl C0=Crbl
xgc_3_25 wwl_3_25 wbl_3_25 rwl_3_25 rbl_3_25 sn_3_25 wos_ros_gc
xrc_wwl_3_25 wwl_3_24 wwl_3_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_25 wbl_2_25 wbl_3_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_25 rwl_3_24 rwl_3_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_25 rbl_2_25 rbl_3_25 rc_unit R0=Rrbl C0=Crbl
xgc_3_26 wwl_3_26 wbl_3_26 rwl_3_26 rbl_3_26 sn_3_26 wos_ros_gc
xrc_wwl_3_26 wwl_3_25 wwl_3_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_26 wbl_2_26 wbl_3_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_26 rwl_3_25 rwl_3_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_26 rbl_2_26 rbl_3_26 rc_unit R0=Rrbl C0=Crbl
xgc_3_27 wwl_3_27 wbl_3_27 rwl_3_27 rbl_3_27 sn_3_27 wos_ros_gc
xrc_wwl_3_27 wwl_3_26 wwl_3_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_27 wbl_2_27 wbl_3_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_27 rwl_3_26 rwl_3_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_27 rbl_2_27 rbl_3_27 rc_unit R0=Rrbl C0=Crbl
xgc_3_28 wwl_3_28 wbl_3_28 rwl_3_28 rbl_3_28 sn_3_28 wos_ros_gc
xrc_wwl_3_28 wwl_3_27 wwl_3_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_28 wbl_2_28 wbl_3_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_28 rwl_3_27 rwl_3_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_28 rbl_2_28 rbl_3_28 rc_unit R0=Rrbl C0=Crbl
xgc_3_29 wwl_3_29 wbl_3_29 rwl_3_29 rbl_3_29 sn_3_29 wos_ros_gc
xrc_wwl_3_29 wwl_3_28 wwl_3_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_29 wbl_2_29 wbl_3_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_29 rwl_3_28 rwl_3_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_29 rbl_2_29 rbl_3_29 rc_unit R0=Rrbl C0=Crbl
xgc_3_30 wwl_3_30 wbl_3_30 rwl_3_30 rbl_3_30 sn_3_30 wos_ros_gc
xrc_wwl_3_30 wwl_3_29 wwl_3_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_30 wbl_2_30 wbl_3_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_30 rwl_3_29 rwl_3_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_30 rbl_2_30 rbl_3_30 rc_unit R0=Rrbl C0=Crbl
xgc_3_31 wwl_3_31 wbl_3_31 rwl_3_31 rbl_3_31 sn_3_31 wos_ros_gc
xrc_wwl_3_31 wwl_3_30 wwl_3_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_3_31 wbl_2_31 wbl_3_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_3_31 rwl_3_30 rwl_3_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_3_31 rbl_2_31 rbl_3_31 rc_unit R0=Rrbl C0=Crbl
xgc_4_0 wwl_4_0 wbl_4_0 rwl_4_0 rbl_4_0 sn_4_0 wos_ros_gc
xrc_wwl_4_0 wwl_4 wwl_4_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_0 wbl_3_0 wbl_4_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_0 rwl_4 rwl_4_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_0 rbl_3_0 rbl_4_0 rc_unit R0=Rrbl C0=Crbl
xgc_4_1 wwl_4_1 wbl_4_1 rwl_4_1 rbl_4_1 sn_4_1 wos_ros_gc
xrc_wwl_4_1 wwl_4_0 wwl_4_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_1 wbl_3_1 wbl_4_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_1 rwl_4_0 rwl_4_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_1 rbl_3_1 rbl_4_1 rc_unit R0=Rrbl C0=Crbl
xgc_4_2 wwl_4_2 wbl_4_2 rwl_4_2 rbl_4_2 sn_4_2 wos_ros_gc
xrc_wwl_4_2 wwl_4_1 wwl_4_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_2 wbl_3_2 wbl_4_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_2 rwl_4_1 rwl_4_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_2 rbl_3_2 rbl_4_2 rc_unit R0=Rrbl C0=Crbl
xgc_4_3 wwl_4_3 wbl_4_3 rwl_4_3 rbl_4_3 sn_4_3 wos_ros_gc
xrc_wwl_4_3 wwl_4_2 wwl_4_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_3 wbl_3_3 wbl_4_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_3 rwl_4_2 rwl_4_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_3 rbl_3_3 rbl_4_3 rc_unit R0=Rrbl C0=Crbl
xgc_4_4 wwl_4_4 wbl_4_4 rwl_4_4 rbl_4_4 sn_4_4 wos_ros_gc
xrc_wwl_4_4 wwl_4_3 wwl_4_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_4 wbl_3_4 wbl_4_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_4 rwl_4_3 rwl_4_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_4 rbl_3_4 rbl_4_4 rc_unit R0=Rrbl C0=Crbl
xgc_4_5 wwl_4_5 wbl_4_5 rwl_4_5 rbl_4_5 sn_4_5 wos_ros_gc
xrc_wwl_4_5 wwl_4_4 wwl_4_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_5 wbl_3_5 wbl_4_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_5 rwl_4_4 rwl_4_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_5 rbl_3_5 rbl_4_5 rc_unit R0=Rrbl C0=Crbl
xgc_4_6 wwl_4_6 wbl_4_6 rwl_4_6 rbl_4_6 sn_4_6 wos_ros_gc
xrc_wwl_4_6 wwl_4_5 wwl_4_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_6 wbl_3_6 wbl_4_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_6 rwl_4_5 rwl_4_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_6 rbl_3_6 rbl_4_6 rc_unit R0=Rrbl C0=Crbl
xgc_4_7 wwl_4_7 wbl_4_7 rwl_4_7 rbl_4_7 sn_4_7 wos_ros_gc
xrc_wwl_4_7 wwl_4_6 wwl_4_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_7 wbl_3_7 wbl_4_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_7 rwl_4_6 rwl_4_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_7 rbl_3_7 rbl_4_7 rc_unit R0=Rrbl C0=Crbl
xgc_4_8 wwl_4_8 wbl_4_8 rwl_4_8 rbl_4_8 sn_4_8 wos_ros_gc
xrc_wwl_4_8 wwl_4_7 wwl_4_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_8 wbl_3_8 wbl_4_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_8 rwl_4_7 rwl_4_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_8 rbl_3_8 rbl_4_8 rc_unit R0=Rrbl C0=Crbl
xgc_4_9 wwl_4_9 wbl_4_9 rwl_4_9 rbl_4_9 sn_4_9 wos_ros_gc
xrc_wwl_4_9 wwl_4_8 wwl_4_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_9 wbl_3_9 wbl_4_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_9 rwl_4_8 rwl_4_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_9 rbl_3_9 rbl_4_9 rc_unit R0=Rrbl C0=Crbl
xgc_4_10 wwl_4_10 wbl_4_10 rwl_4_10 rbl_4_10 sn_4_10 wos_ros_gc
xrc_wwl_4_10 wwl_4_9 wwl_4_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_10 wbl_3_10 wbl_4_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_10 rwl_4_9 rwl_4_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_10 rbl_3_10 rbl_4_10 rc_unit R0=Rrbl C0=Crbl
xgc_4_11 wwl_4_11 wbl_4_11 rwl_4_11 rbl_4_11 sn_4_11 wos_ros_gc
xrc_wwl_4_11 wwl_4_10 wwl_4_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_11 wbl_3_11 wbl_4_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_11 rwl_4_10 rwl_4_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_11 rbl_3_11 rbl_4_11 rc_unit R0=Rrbl C0=Crbl
xgc_4_12 wwl_4_12 wbl_4_12 rwl_4_12 rbl_4_12 sn_4_12 wos_ros_gc
xrc_wwl_4_12 wwl_4_11 wwl_4_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_12 wbl_3_12 wbl_4_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_12 rwl_4_11 rwl_4_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_12 rbl_3_12 rbl_4_12 rc_unit R0=Rrbl C0=Crbl
xgc_4_13 wwl_4_13 wbl_4_13 rwl_4_13 rbl_4_13 sn_4_13 wos_ros_gc
xrc_wwl_4_13 wwl_4_12 wwl_4_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_13 wbl_3_13 wbl_4_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_13 rwl_4_12 rwl_4_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_13 rbl_3_13 rbl_4_13 rc_unit R0=Rrbl C0=Crbl
xgc_4_14 wwl_4_14 wbl_4_14 rwl_4_14 rbl_4_14 sn_4_14 wos_ros_gc
xrc_wwl_4_14 wwl_4_13 wwl_4_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_14 wbl_3_14 wbl_4_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_14 rwl_4_13 rwl_4_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_14 rbl_3_14 rbl_4_14 rc_unit R0=Rrbl C0=Crbl
xgc_4_15 wwl_4_15 wbl_4_15 rwl_4_15 rbl_4_15 sn_4_15 wos_ros_gc
xrc_wwl_4_15 wwl_4_14 wwl_4_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_15 wbl_3_15 wbl_4_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_15 rwl_4_14 rwl_4_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_15 rbl_3_15 rbl_4_15 rc_unit R0=Rrbl C0=Crbl
xgc_4_16 wwl_4_16 wbl_4_16 rwl_4_16 rbl_4_16 sn_4_16 wos_ros_gc
xrc_wwl_4_16 wwl_4_15 wwl_4_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_16 wbl_3_16 wbl_4_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_16 rwl_4_15 rwl_4_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_16 rbl_3_16 rbl_4_16 rc_unit R0=Rrbl C0=Crbl
xgc_4_17 wwl_4_17 wbl_4_17 rwl_4_17 rbl_4_17 sn_4_17 wos_ros_gc
xrc_wwl_4_17 wwl_4_16 wwl_4_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_17 wbl_3_17 wbl_4_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_17 rwl_4_16 rwl_4_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_17 rbl_3_17 rbl_4_17 rc_unit R0=Rrbl C0=Crbl
xgc_4_18 wwl_4_18 wbl_4_18 rwl_4_18 rbl_4_18 sn_4_18 wos_ros_gc
xrc_wwl_4_18 wwl_4_17 wwl_4_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_18 wbl_3_18 wbl_4_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_18 rwl_4_17 rwl_4_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_18 rbl_3_18 rbl_4_18 rc_unit R0=Rrbl C0=Crbl
xgc_4_19 wwl_4_19 wbl_4_19 rwl_4_19 rbl_4_19 sn_4_19 wos_ros_gc
xrc_wwl_4_19 wwl_4_18 wwl_4_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_19 wbl_3_19 wbl_4_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_19 rwl_4_18 rwl_4_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_19 rbl_3_19 rbl_4_19 rc_unit R0=Rrbl C0=Crbl
xgc_4_20 wwl_4_20 wbl_4_20 rwl_4_20 rbl_4_20 sn_4_20 wos_ros_gc
xrc_wwl_4_20 wwl_4_19 wwl_4_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_20 wbl_3_20 wbl_4_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_20 rwl_4_19 rwl_4_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_20 rbl_3_20 rbl_4_20 rc_unit R0=Rrbl C0=Crbl
xgc_4_21 wwl_4_21 wbl_4_21 rwl_4_21 rbl_4_21 sn_4_21 wos_ros_gc
xrc_wwl_4_21 wwl_4_20 wwl_4_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_21 wbl_3_21 wbl_4_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_21 rwl_4_20 rwl_4_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_21 rbl_3_21 rbl_4_21 rc_unit R0=Rrbl C0=Crbl
xgc_4_22 wwl_4_22 wbl_4_22 rwl_4_22 rbl_4_22 sn_4_22 wos_ros_gc
xrc_wwl_4_22 wwl_4_21 wwl_4_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_22 wbl_3_22 wbl_4_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_22 rwl_4_21 rwl_4_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_22 rbl_3_22 rbl_4_22 rc_unit R0=Rrbl C0=Crbl
xgc_4_23 wwl_4_23 wbl_4_23 rwl_4_23 rbl_4_23 sn_4_23 wos_ros_gc
xrc_wwl_4_23 wwl_4_22 wwl_4_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_23 wbl_3_23 wbl_4_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_23 rwl_4_22 rwl_4_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_23 rbl_3_23 rbl_4_23 rc_unit R0=Rrbl C0=Crbl
xgc_4_24 wwl_4_24 wbl_4_24 rwl_4_24 rbl_4_24 sn_4_24 wos_ros_gc
xrc_wwl_4_24 wwl_4_23 wwl_4_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_24 wbl_3_24 wbl_4_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_24 rwl_4_23 rwl_4_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_24 rbl_3_24 rbl_4_24 rc_unit R0=Rrbl C0=Crbl
xgc_4_25 wwl_4_25 wbl_4_25 rwl_4_25 rbl_4_25 sn_4_25 wos_ros_gc
xrc_wwl_4_25 wwl_4_24 wwl_4_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_25 wbl_3_25 wbl_4_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_25 rwl_4_24 rwl_4_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_25 rbl_3_25 rbl_4_25 rc_unit R0=Rrbl C0=Crbl
xgc_4_26 wwl_4_26 wbl_4_26 rwl_4_26 rbl_4_26 sn_4_26 wos_ros_gc
xrc_wwl_4_26 wwl_4_25 wwl_4_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_26 wbl_3_26 wbl_4_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_26 rwl_4_25 rwl_4_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_26 rbl_3_26 rbl_4_26 rc_unit R0=Rrbl C0=Crbl
xgc_4_27 wwl_4_27 wbl_4_27 rwl_4_27 rbl_4_27 sn_4_27 wos_ros_gc
xrc_wwl_4_27 wwl_4_26 wwl_4_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_27 wbl_3_27 wbl_4_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_27 rwl_4_26 rwl_4_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_27 rbl_3_27 rbl_4_27 rc_unit R0=Rrbl C0=Crbl
xgc_4_28 wwl_4_28 wbl_4_28 rwl_4_28 rbl_4_28 sn_4_28 wos_ros_gc
xrc_wwl_4_28 wwl_4_27 wwl_4_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_28 wbl_3_28 wbl_4_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_28 rwl_4_27 rwl_4_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_28 rbl_3_28 rbl_4_28 rc_unit R0=Rrbl C0=Crbl
xgc_4_29 wwl_4_29 wbl_4_29 rwl_4_29 rbl_4_29 sn_4_29 wos_ros_gc
xrc_wwl_4_29 wwl_4_28 wwl_4_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_29 wbl_3_29 wbl_4_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_29 rwl_4_28 rwl_4_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_29 rbl_3_29 rbl_4_29 rc_unit R0=Rrbl C0=Crbl
xgc_4_30 wwl_4_30 wbl_4_30 rwl_4_30 rbl_4_30 sn_4_30 wos_ros_gc
xrc_wwl_4_30 wwl_4_29 wwl_4_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_30 wbl_3_30 wbl_4_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_30 rwl_4_29 rwl_4_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_30 rbl_3_30 rbl_4_30 rc_unit R0=Rrbl C0=Crbl
xgc_4_31 wwl_4_31 wbl_4_31 rwl_4_31 rbl_4_31 sn_4_31 wos_ros_gc
xrc_wwl_4_31 wwl_4_30 wwl_4_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_4_31 wbl_3_31 wbl_4_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_4_31 rwl_4_30 rwl_4_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_4_31 rbl_3_31 rbl_4_31 rc_unit R0=Rrbl C0=Crbl
xgc_5_0 wwl_5_0 wbl_5_0 rwl_5_0 rbl_5_0 sn_5_0 wos_ros_gc
xrc_wwl_5_0 wwl_5 wwl_5_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_0 wbl_4_0 wbl_5_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_0 rwl_5 rwl_5_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_0 rbl_4_0 rbl_5_0 rc_unit R0=Rrbl C0=Crbl
xgc_5_1 wwl_5_1 wbl_5_1 rwl_5_1 rbl_5_1 sn_5_1 wos_ros_gc
xrc_wwl_5_1 wwl_5_0 wwl_5_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_1 wbl_4_1 wbl_5_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_1 rwl_5_0 rwl_5_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_1 rbl_4_1 rbl_5_1 rc_unit R0=Rrbl C0=Crbl
xgc_5_2 wwl_5_2 wbl_5_2 rwl_5_2 rbl_5_2 sn_5_2 wos_ros_gc
xrc_wwl_5_2 wwl_5_1 wwl_5_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_2 wbl_4_2 wbl_5_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_2 rwl_5_1 rwl_5_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_2 rbl_4_2 rbl_5_2 rc_unit R0=Rrbl C0=Crbl
xgc_5_3 wwl_5_3 wbl_5_3 rwl_5_3 rbl_5_3 sn_5_3 wos_ros_gc
xrc_wwl_5_3 wwl_5_2 wwl_5_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_3 wbl_4_3 wbl_5_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_3 rwl_5_2 rwl_5_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_3 rbl_4_3 rbl_5_3 rc_unit R0=Rrbl C0=Crbl
xgc_5_4 wwl_5_4 wbl_5_4 rwl_5_4 rbl_5_4 sn_5_4 wos_ros_gc
xrc_wwl_5_4 wwl_5_3 wwl_5_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_4 wbl_4_4 wbl_5_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_4 rwl_5_3 rwl_5_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_4 rbl_4_4 rbl_5_4 rc_unit R0=Rrbl C0=Crbl
xgc_5_5 wwl_5_5 wbl_5_5 rwl_5_5 rbl_5_5 sn_5_5 wos_ros_gc
xrc_wwl_5_5 wwl_5_4 wwl_5_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_5 wbl_4_5 wbl_5_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_5 rwl_5_4 rwl_5_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_5 rbl_4_5 rbl_5_5 rc_unit R0=Rrbl C0=Crbl
xgc_5_6 wwl_5_6 wbl_5_6 rwl_5_6 rbl_5_6 sn_5_6 wos_ros_gc
xrc_wwl_5_6 wwl_5_5 wwl_5_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_6 wbl_4_6 wbl_5_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_6 rwl_5_5 rwl_5_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_6 rbl_4_6 rbl_5_6 rc_unit R0=Rrbl C0=Crbl
xgc_5_7 wwl_5_7 wbl_5_7 rwl_5_7 rbl_5_7 sn_5_7 wos_ros_gc
xrc_wwl_5_7 wwl_5_6 wwl_5_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_7 wbl_4_7 wbl_5_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_7 rwl_5_6 rwl_5_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_7 rbl_4_7 rbl_5_7 rc_unit R0=Rrbl C0=Crbl
xgc_5_8 wwl_5_8 wbl_5_8 rwl_5_8 rbl_5_8 sn_5_8 wos_ros_gc
xrc_wwl_5_8 wwl_5_7 wwl_5_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_8 wbl_4_8 wbl_5_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_8 rwl_5_7 rwl_5_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_8 rbl_4_8 rbl_5_8 rc_unit R0=Rrbl C0=Crbl
xgc_5_9 wwl_5_9 wbl_5_9 rwl_5_9 rbl_5_9 sn_5_9 wos_ros_gc
xrc_wwl_5_9 wwl_5_8 wwl_5_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_9 wbl_4_9 wbl_5_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_9 rwl_5_8 rwl_5_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_9 rbl_4_9 rbl_5_9 rc_unit R0=Rrbl C0=Crbl
xgc_5_10 wwl_5_10 wbl_5_10 rwl_5_10 rbl_5_10 sn_5_10 wos_ros_gc
xrc_wwl_5_10 wwl_5_9 wwl_5_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_10 wbl_4_10 wbl_5_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_10 rwl_5_9 rwl_5_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_10 rbl_4_10 rbl_5_10 rc_unit R0=Rrbl C0=Crbl
xgc_5_11 wwl_5_11 wbl_5_11 rwl_5_11 rbl_5_11 sn_5_11 wos_ros_gc
xrc_wwl_5_11 wwl_5_10 wwl_5_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_11 wbl_4_11 wbl_5_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_11 rwl_5_10 rwl_5_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_11 rbl_4_11 rbl_5_11 rc_unit R0=Rrbl C0=Crbl
xgc_5_12 wwl_5_12 wbl_5_12 rwl_5_12 rbl_5_12 sn_5_12 wos_ros_gc
xrc_wwl_5_12 wwl_5_11 wwl_5_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_12 wbl_4_12 wbl_5_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_12 rwl_5_11 rwl_5_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_12 rbl_4_12 rbl_5_12 rc_unit R0=Rrbl C0=Crbl
xgc_5_13 wwl_5_13 wbl_5_13 rwl_5_13 rbl_5_13 sn_5_13 wos_ros_gc
xrc_wwl_5_13 wwl_5_12 wwl_5_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_13 wbl_4_13 wbl_5_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_13 rwl_5_12 rwl_5_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_13 rbl_4_13 rbl_5_13 rc_unit R0=Rrbl C0=Crbl
xgc_5_14 wwl_5_14 wbl_5_14 rwl_5_14 rbl_5_14 sn_5_14 wos_ros_gc
xrc_wwl_5_14 wwl_5_13 wwl_5_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_14 wbl_4_14 wbl_5_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_14 rwl_5_13 rwl_5_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_14 rbl_4_14 rbl_5_14 rc_unit R0=Rrbl C0=Crbl
xgc_5_15 wwl_5_15 wbl_5_15 rwl_5_15 rbl_5_15 sn_5_15 wos_ros_gc
xrc_wwl_5_15 wwl_5_14 wwl_5_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_15 wbl_4_15 wbl_5_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_15 rwl_5_14 rwl_5_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_15 rbl_4_15 rbl_5_15 rc_unit R0=Rrbl C0=Crbl
xgc_5_16 wwl_5_16 wbl_5_16 rwl_5_16 rbl_5_16 sn_5_16 wos_ros_gc
xrc_wwl_5_16 wwl_5_15 wwl_5_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_16 wbl_4_16 wbl_5_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_16 rwl_5_15 rwl_5_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_16 rbl_4_16 rbl_5_16 rc_unit R0=Rrbl C0=Crbl
xgc_5_17 wwl_5_17 wbl_5_17 rwl_5_17 rbl_5_17 sn_5_17 wos_ros_gc
xrc_wwl_5_17 wwl_5_16 wwl_5_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_17 wbl_4_17 wbl_5_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_17 rwl_5_16 rwl_5_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_17 rbl_4_17 rbl_5_17 rc_unit R0=Rrbl C0=Crbl
xgc_5_18 wwl_5_18 wbl_5_18 rwl_5_18 rbl_5_18 sn_5_18 wos_ros_gc
xrc_wwl_5_18 wwl_5_17 wwl_5_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_18 wbl_4_18 wbl_5_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_18 rwl_5_17 rwl_5_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_18 rbl_4_18 rbl_5_18 rc_unit R0=Rrbl C0=Crbl
xgc_5_19 wwl_5_19 wbl_5_19 rwl_5_19 rbl_5_19 sn_5_19 wos_ros_gc
xrc_wwl_5_19 wwl_5_18 wwl_5_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_19 wbl_4_19 wbl_5_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_19 rwl_5_18 rwl_5_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_19 rbl_4_19 rbl_5_19 rc_unit R0=Rrbl C0=Crbl
xgc_5_20 wwl_5_20 wbl_5_20 rwl_5_20 rbl_5_20 sn_5_20 wos_ros_gc
xrc_wwl_5_20 wwl_5_19 wwl_5_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_20 wbl_4_20 wbl_5_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_20 rwl_5_19 rwl_5_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_20 rbl_4_20 rbl_5_20 rc_unit R0=Rrbl C0=Crbl
xgc_5_21 wwl_5_21 wbl_5_21 rwl_5_21 rbl_5_21 sn_5_21 wos_ros_gc
xrc_wwl_5_21 wwl_5_20 wwl_5_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_21 wbl_4_21 wbl_5_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_21 rwl_5_20 rwl_5_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_21 rbl_4_21 rbl_5_21 rc_unit R0=Rrbl C0=Crbl
xgc_5_22 wwl_5_22 wbl_5_22 rwl_5_22 rbl_5_22 sn_5_22 wos_ros_gc
xrc_wwl_5_22 wwl_5_21 wwl_5_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_22 wbl_4_22 wbl_5_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_22 rwl_5_21 rwl_5_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_22 rbl_4_22 rbl_5_22 rc_unit R0=Rrbl C0=Crbl
xgc_5_23 wwl_5_23 wbl_5_23 rwl_5_23 rbl_5_23 sn_5_23 wos_ros_gc
xrc_wwl_5_23 wwl_5_22 wwl_5_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_23 wbl_4_23 wbl_5_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_23 rwl_5_22 rwl_5_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_23 rbl_4_23 rbl_5_23 rc_unit R0=Rrbl C0=Crbl
xgc_5_24 wwl_5_24 wbl_5_24 rwl_5_24 rbl_5_24 sn_5_24 wos_ros_gc
xrc_wwl_5_24 wwl_5_23 wwl_5_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_24 wbl_4_24 wbl_5_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_24 rwl_5_23 rwl_5_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_24 rbl_4_24 rbl_5_24 rc_unit R0=Rrbl C0=Crbl
xgc_5_25 wwl_5_25 wbl_5_25 rwl_5_25 rbl_5_25 sn_5_25 wos_ros_gc
xrc_wwl_5_25 wwl_5_24 wwl_5_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_25 wbl_4_25 wbl_5_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_25 rwl_5_24 rwl_5_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_25 rbl_4_25 rbl_5_25 rc_unit R0=Rrbl C0=Crbl
xgc_5_26 wwl_5_26 wbl_5_26 rwl_5_26 rbl_5_26 sn_5_26 wos_ros_gc
xrc_wwl_5_26 wwl_5_25 wwl_5_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_26 wbl_4_26 wbl_5_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_26 rwl_5_25 rwl_5_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_26 rbl_4_26 rbl_5_26 rc_unit R0=Rrbl C0=Crbl
xgc_5_27 wwl_5_27 wbl_5_27 rwl_5_27 rbl_5_27 sn_5_27 wos_ros_gc
xrc_wwl_5_27 wwl_5_26 wwl_5_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_27 wbl_4_27 wbl_5_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_27 rwl_5_26 rwl_5_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_27 rbl_4_27 rbl_5_27 rc_unit R0=Rrbl C0=Crbl
xgc_5_28 wwl_5_28 wbl_5_28 rwl_5_28 rbl_5_28 sn_5_28 wos_ros_gc
xrc_wwl_5_28 wwl_5_27 wwl_5_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_28 wbl_4_28 wbl_5_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_28 rwl_5_27 rwl_5_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_28 rbl_4_28 rbl_5_28 rc_unit R0=Rrbl C0=Crbl
xgc_5_29 wwl_5_29 wbl_5_29 rwl_5_29 rbl_5_29 sn_5_29 wos_ros_gc
xrc_wwl_5_29 wwl_5_28 wwl_5_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_29 wbl_4_29 wbl_5_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_29 rwl_5_28 rwl_5_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_29 rbl_4_29 rbl_5_29 rc_unit R0=Rrbl C0=Crbl
xgc_5_30 wwl_5_30 wbl_5_30 rwl_5_30 rbl_5_30 sn_5_30 wos_ros_gc
xrc_wwl_5_30 wwl_5_29 wwl_5_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_30 wbl_4_30 wbl_5_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_30 rwl_5_29 rwl_5_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_30 rbl_4_30 rbl_5_30 rc_unit R0=Rrbl C0=Crbl
xgc_5_31 wwl_5_31 wbl_5_31 rwl_5_31 rbl_5_31 sn_5_31 wos_ros_gc
xrc_wwl_5_31 wwl_5_30 wwl_5_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_5_31 wbl_4_31 wbl_5_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_5_31 rwl_5_30 rwl_5_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_5_31 rbl_4_31 rbl_5_31 rc_unit R0=Rrbl C0=Crbl
xgc_6_0 wwl_6_0 wbl_6_0 rwl_6_0 rbl_6_0 sn_6_0 wos_ros_gc
xrc_wwl_6_0 wwl_6 wwl_6_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_0 wbl_5_0 wbl_6_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_0 rwl_6 rwl_6_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_0 rbl_5_0 rbl_6_0 rc_unit R0=Rrbl C0=Crbl
xgc_6_1 wwl_6_1 wbl_6_1 rwl_6_1 rbl_6_1 sn_6_1 wos_ros_gc
xrc_wwl_6_1 wwl_6_0 wwl_6_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_1 wbl_5_1 wbl_6_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_1 rwl_6_0 rwl_6_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_1 rbl_5_1 rbl_6_1 rc_unit R0=Rrbl C0=Crbl
xgc_6_2 wwl_6_2 wbl_6_2 rwl_6_2 rbl_6_2 sn_6_2 wos_ros_gc
xrc_wwl_6_2 wwl_6_1 wwl_6_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_2 wbl_5_2 wbl_6_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_2 rwl_6_1 rwl_6_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_2 rbl_5_2 rbl_6_2 rc_unit R0=Rrbl C0=Crbl
xgc_6_3 wwl_6_3 wbl_6_3 rwl_6_3 rbl_6_3 sn_6_3 wos_ros_gc
xrc_wwl_6_3 wwl_6_2 wwl_6_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_3 wbl_5_3 wbl_6_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_3 rwl_6_2 rwl_6_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_3 rbl_5_3 rbl_6_3 rc_unit R0=Rrbl C0=Crbl
xgc_6_4 wwl_6_4 wbl_6_4 rwl_6_4 rbl_6_4 sn_6_4 wos_ros_gc
xrc_wwl_6_4 wwl_6_3 wwl_6_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_4 wbl_5_4 wbl_6_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_4 rwl_6_3 rwl_6_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_4 rbl_5_4 rbl_6_4 rc_unit R0=Rrbl C0=Crbl
xgc_6_5 wwl_6_5 wbl_6_5 rwl_6_5 rbl_6_5 sn_6_5 wos_ros_gc
xrc_wwl_6_5 wwl_6_4 wwl_6_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_5 wbl_5_5 wbl_6_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_5 rwl_6_4 rwl_6_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_5 rbl_5_5 rbl_6_5 rc_unit R0=Rrbl C0=Crbl
xgc_6_6 wwl_6_6 wbl_6_6 rwl_6_6 rbl_6_6 sn_6_6 wos_ros_gc
xrc_wwl_6_6 wwl_6_5 wwl_6_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_6 wbl_5_6 wbl_6_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_6 rwl_6_5 rwl_6_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_6 rbl_5_6 rbl_6_6 rc_unit R0=Rrbl C0=Crbl
xgc_6_7 wwl_6_7 wbl_6_7 rwl_6_7 rbl_6_7 sn_6_7 wos_ros_gc
xrc_wwl_6_7 wwl_6_6 wwl_6_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_7 wbl_5_7 wbl_6_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_7 rwl_6_6 rwl_6_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_7 rbl_5_7 rbl_6_7 rc_unit R0=Rrbl C0=Crbl
xgc_6_8 wwl_6_8 wbl_6_8 rwl_6_8 rbl_6_8 sn_6_8 wos_ros_gc
xrc_wwl_6_8 wwl_6_7 wwl_6_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_8 wbl_5_8 wbl_6_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_8 rwl_6_7 rwl_6_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_8 rbl_5_8 rbl_6_8 rc_unit R0=Rrbl C0=Crbl
xgc_6_9 wwl_6_9 wbl_6_9 rwl_6_9 rbl_6_9 sn_6_9 wos_ros_gc
xrc_wwl_6_9 wwl_6_8 wwl_6_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_9 wbl_5_9 wbl_6_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_9 rwl_6_8 rwl_6_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_9 rbl_5_9 rbl_6_9 rc_unit R0=Rrbl C0=Crbl
xgc_6_10 wwl_6_10 wbl_6_10 rwl_6_10 rbl_6_10 sn_6_10 wos_ros_gc
xrc_wwl_6_10 wwl_6_9 wwl_6_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_10 wbl_5_10 wbl_6_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_10 rwl_6_9 rwl_6_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_10 rbl_5_10 rbl_6_10 rc_unit R0=Rrbl C0=Crbl
xgc_6_11 wwl_6_11 wbl_6_11 rwl_6_11 rbl_6_11 sn_6_11 wos_ros_gc
xrc_wwl_6_11 wwl_6_10 wwl_6_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_11 wbl_5_11 wbl_6_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_11 rwl_6_10 rwl_6_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_11 rbl_5_11 rbl_6_11 rc_unit R0=Rrbl C0=Crbl
xgc_6_12 wwl_6_12 wbl_6_12 rwl_6_12 rbl_6_12 sn_6_12 wos_ros_gc
xrc_wwl_6_12 wwl_6_11 wwl_6_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_12 wbl_5_12 wbl_6_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_12 rwl_6_11 rwl_6_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_12 rbl_5_12 rbl_6_12 rc_unit R0=Rrbl C0=Crbl
xgc_6_13 wwl_6_13 wbl_6_13 rwl_6_13 rbl_6_13 sn_6_13 wos_ros_gc
xrc_wwl_6_13 wwl_6_12 wwl_6_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_13 wbl_5_13 wbl_6_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_13 rwl_6_12 rwl_6_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_13 rbl_5_13 rbl_6_13 rc_unit R0=Rrbl C0=Crbl
xgc_6_14 wwl_6_14 wbl_6_14 rwl_6_14 rbl_6_14 sn_6_14 wos_ros_gc
xrc_wwl_6_14 wwl_6_13 wwl_6_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_14 wbl_5_14 wbl_6_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_14 rwl_6_13 rwl_6_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_14 rbl_5_14 rbl_6_14 rc_unit R0=Rrbl C0=Crbl
xgc_6_15 wwl_6_15 wbl_6_15 rwl_6_15 rbl_6_15 sn_6_15 wos_ros_gc
xrc_wwl_6_15 wwl_6_14 wwl_6_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_15 wbl_5_15 wbl_6_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_15 rwl_6_14 rwl_6_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_15 rbl_5_15 rbl_6_15 rc_unit R0=Rrbl C0=Crbl
xgc_6_16 wwl_6_16 wbl_6_16 rwl_6_16 rbl_6_16 sn_6_16 wos_ros_gc
xrc_wwl_6_16 wwl_6_15 wwl_6_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_16 wbl_5_16 wbl_6_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_16 rwl_6_15 rwl_6_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_16 rbl_5_16 rbl_6_16 rc_unit R0=Rrbl C0=Crbl
xgc_6_17 wwl_6_17 wbl_6_17 rwl_6_17 rbl_6_17 sn_6_17 wos_ros_gc
xrc_wwl_6_17 wwl_6_16 wwl_6_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_17 wbl_5_17 wbl_6_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_17 rwl_6_16 rwl_6_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_17 rbl_5_17 rbl_6_17 rc_unit R0=Rrbl C0=Crbl
xgc_6_18 wwl_6_18 wbl_6_18 rwl_6_18 rbl_6_18 sn_6_18 wos_ros_gc
xrc_wwl_6_18 wwl_6_17 wwl_6_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_18 wbl_5_18 wbl_6_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_18 rwl_6_17 rwl_6_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_18 rbl_5_18 rbl_6_18 rc_unit R0=Rrbl C0=Crbl
xgc_6_19 wwl_6_19 wbl_6_19 rwl_6_19 rbl_6_19 sn_6_19 wos_ros_gc
xrc_wwl_6_19 wwl_6_18 wwl_6_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_19 wbl_5_19 wbl_6_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_19 rwl_6_18 rwl_6_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_19 rbl_5_19 rbl_6_19 rc_unit R0=Rrbl C0=Crbl
xgc_6_20 wwl_6_20 wbl_6_20 rwl_6_20 rbl_6_20 sn_6_20 wos_ros_gc
xrc_wwl_6_20 wwl_6_19 wwl_6_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_20 wbl_5_20 wbl_6_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_20 rwl_6_19 rwl_6_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_20 rbl_5_20 rbl_6_20 rc_unit R0=Rrbl C0=Crbl
xgc_6_21 wwl_6_21 wbl_6_21 rwl_6_21 rbl_6_21 sn_6_21 wos_ros_gc
xrc_wwl_6_21 wwl_6_20 wwl_6_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_21 wbl_5_21 wbl_6_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_21 rwl_6_20 rwl_6_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_21 rbl_5_21 rbl_6_21 rc_unit R0=Rrbl C0=Crbl
xgc_6_22 wwl_6_22 wbl_6_22 rwl_6_22 rbl_6_22 sn_6_22 wos_ros_gc
xrc_wwl_6_22 wwl_6_21 wwl_6_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_22 wbl_5_22 wbl_6_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_22 rwl_6_21 rwl_6_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_22 rbl_5_22 rbl_6_22 rc_unit R0=Rrbl C0=Crbl
xgc_6_23 wwl_6_23 wbl_6_23 rwl_6_23 rbl_6_23 sn_6_23 wos_ros_gc
xrc_wwl_6_23 wwl_6_22 wwl_6_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_23 wbl_5_23 wbl_6_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_23 rwl_6_22 rwl_6_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_23 rbl_5_23 rbl_6_23 rc_unit R0=Rrbl C0=Crbl
xgc_6_24 wwl_6_24 wbl_6_24 rwl_6_24 rbl_6_24 sn_6_24 wos_ros_gc
xrc_wwl_6_24 wwl_6_23 wwl_6_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_24 wbl_5_24 wbl_6_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_24 rwl_6_23 rwl_6_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_24 rbl_5_24 rbl_6_24 rc_unit R0=Rrbl C0=Crbl
xgc_6_25 wwl_6_25 wbl_6_25 rwl_6_25 rbl_6_25 sn_6_25 wos_ros_gc
xrc_wwl_6_25 wwl_6_24 wwl_6_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_25 wbl_5_25 wbl_6_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_25 rwl_6_24 rwl_6_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_25 rbl_5_25 rbl_6_25 rc_unit R0=Rrbl C0=Crbl
xgc_6_26 wwl_6_26 wbl_6_26 rwl_6_26 rbl_6_26 sn_6_26 wos_ros_gc
xrc_wwl_6_26 wwl_6_25 wwl_6_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_26 wbl_5_26 wbl_6_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_26 rwl_6_25 rwl_6_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_26 rbl_5_26 rbl_6_26 rc_unit R0=Rrbl C0=Crbl
xgc_6_27 wwl_6_27 wbl_6_27 rwl_6_27 rbl_6_27 sn_6_27 wos_ros_gc
xrc_wwl_6_27 wwl_6_26 wwl_6_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_27 wbl_5_27 wbl_6_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_27 rwl_6_26 rwl_6_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_27 rbl_5_27 rbl_6_27 rc_unit R0=Rrbl C0=Crbl
xgc_6_28 wwl_6_28 wbl_6_28 rwl_6_28 rbl_6_28 sn_6_28 wos_ros_gc
xrc_wwl_6_28 wwl_6_27 wwl_6_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_28 wbl_5_28 wbl_6_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_28 rwl_6_27 rwl_6_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_28 rbl_5_28 rbl_6_28 rc_unit R0=Rrbl C0=Crbl
xgc_6_29 wwl_6_29 wbl_6_29 rwl_6_29 rbl_6_29 sn_6_29 wos_ros_gc
xrc_wwl_6_29 wwl_6_28 wwl_6_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_29 wbl_5_29 wbl_6_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_29 rwl_6_28 rwl_6_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_29 rbl_5_29 rbl_6_29 rc_unit R0=Rrbl C0=Crbl
xgc_6_30 wwl_6_30 wbl_6_30 rwl_6_30 rbl_6_30 sn_6_30 wos_ros_gc
xrc_wwl_6_30 wwl_6_29 wwl_6_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_30 wbl_5_30 wbl_6_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_30 rwl_6_29 rwl_6_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_30 rbl_5_30 rbl_6_30 rc_unit R0=Rrbl C0=Crbl
xgc_6_31 wwl_6_31 wbl_6_31 rwl_6_31 rbl_6_31 sn_6_31 wos_ros_gc
xrc_wwl_6_31 wwl_6_30 wwl_6_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_6_31 wbl_5_31 wbl_6_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_6_31 rwl_6_30 rwl_6_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_6_31 rbl_5_31 rbl_6_31 rc_unit R0=Rrbl C0=Crbl
xgc_7_0 wwl_7_0 wbl_7_0 rwl_7_0 rbl_7_0 sn_7_0 wos_ros_gc
xrc_wwl_7_0 wwl_7 wwl_7_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_0 wbl_6_0 wbl_7_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_0 rwl_7 rwl_7_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_0 rbl_6_0 rbl_7_0 rc_unit R0=Rrbl C0=Crbl
xgc_7_1 wwl_7_1 wbl_7_1 rwl_7_1 rbl_7_1 sn_7_1 wos_ros_gc
xrc_wwl_7_1 wwl_7_0 wwl_7_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_1 wbl_6_1 wbl_7_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_1 rwl_7_0 rwl_7_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_1 rbl_6_1 rbl_7_1 rc_unit R0=Rrbl C0=Crbl
xgc_7_2 wwl_7_2 wbl_7_2 rwl_7_2 rbl_7_2 sn_7_2 wos_ros_gc
xrc_wwl_7_2 wwl_7_1 wwl_7_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_2 wbl_6_2 wbl_7_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_2 rwl_7_1 rwl_7_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_2 rbl_6_2 rbl_7_2 rc_unit R0=Rrbl C0=Crbl
xgc_7_3 wwl_7_3 wbl_7_3 rwl_7_3 rbl_7_3 sn_7_3 wos_ros_gc
xrc_wwl_7_3 wwl_7_2 wwl_7_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_3 wbl_6_3 wbl_7_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_3 rwl_7_2 rwl_7_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_3 rbl_6_3 rbl_7_3 rc_unit R0=Rrbl C0=Crbl
xgc_7_4 wwl_7_4 wbl_7_4 rwl_7_4 rbl_7_4 sn_7_4 wos_ros_gc
xrc_wwl_7_4 wwl_7_3 wwl_7_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_4 wbl_6_4 wbl_7_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_4 rwl_7_3 rwl_7_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_4 rbl_6_4 rbl_7_4 rc_unit R0=Rrbl C0=Crbl
xgc_7_5 wwl_7_5 wbl_7_5 rwl_7_5 rbl_7_5 sn_7_5 wos_ros_gc
xrc_wwl_7_5 wwl_7_4 wwl_7_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_5 wbl_6_5 wbl_7_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_5 rwl_7_4 rwl_7_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_5 rbl_6_5 rbl_7_5 rc_unit R0=Rrbl C0=Crbl
xgc_7_6 wwl_7_6 wbl_7_6 rwl_7_6 rbl_7_6 sn_7_6 wos_ros_gc
xrc_wwl_7_6 wwl_7_5 wwl_7_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_6 wbl_6_6 wbl_7_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_6 rwl_7_5 rwl_7_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_6 rbl_6_6 rbl_7_6 rc_unit R0=Rrbl C0=Crbl
xgc_7_7 wwl_7_7 wbl_7_7 rwl_7_7 rbl_7_7 sn_7_7 wos_ros_gc
xrc_wwl_7_7 wwl_7_6 wwl_7_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_7 wbl_6_7 wbl_7_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_7 rwl_7_6 rwl_7_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_7 rbl_6_7 rbl_7_7 rc_unit R0=Rrbl C0=Crbl
xgc_7_8 wwl_7_8 wbl_7_8 rwl_7_8 rbl_7_8 sn_7_8 wos_ros_gc
xrc_wwl_7_8 wwl_7_7 wwl_7_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_8 wbl_6_8 wbl_7_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_8 rwl_7_7 rwl_7_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_8 rbl_6_8 rbl_7_8 rc_unit R0=Rrbl C0=Crbl
xgc_7_9 wwl_7_9 wbl_7_9 rwl_7_9 rbl_7_9 sn_7_9 wos_ros_gc
xrc_wwl_7_9 wwl_7_8 wwl_7_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_9 wbl_6_9 wbl_7_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_9 rwl_7_8 rwl_7_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_9 rbl_6_9 rbl_7_9 rc_unit R0=Rrbl C0=Crbl
xgc_7_10 wwl_7_10 wbl_7_10 rwl_7_10 rbl_7_10 sn_7_10 wos_ros_gc
xrc_wwl_7_10 wwl_7_9 wwl_7_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_10 wbl_6_10 wbl_7_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_10 rwl_7_9 rwl_7_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_10 rbl_6_10 rbl_7_10 rc_unit R0=Rrbl C0=Crbl
xgc_7_11 wwl_7_11 wbl_7_11 rwl_7_11 rbl_7_11 sn_7_11 wos_ros_gc
xrc_wwl_7_11 wwl_7_10 wwl_7_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_11 wbl_6_11 wbl_7_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_11 rwl_7_10 rwl_7_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_11 rbl_6_11 rbl_7_11 rc_unit R0=Rrbl C0=Crbl
xgc_7_12 wwl_7_12 wbl_7_12 rwl_7_12 rbl_7_12 sn_7_12 wos_ros_gc
xrc_wwl_7_12 wwl_7_11 wwl_7_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_12 wbl_6_12 wbl_7_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_12 rwl_7_11 rwl_7_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_12 rbl_6_12 rbl_7_12 rc_unit R0=Rrbl C0=Crbl
xgc_7_13 wwl_7_13 wbl_7_13 rwl_7_13 rbl_7_13 sn_7_13 wos_ros_gc
xrc_wwl_7_13 wwl_7_12 wwl_7_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_13 wbl_6_13 wbl_7_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_13 rwl_7_12 rwl_7_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_13 rbl_6_13 rbl_7_13 rc_unit R0=Rrbl C0=Crbl
xgc_7_14 wwl_7_14 wbl_7_14 rwl_7_14 rbl_7_14 sn_7_14 wos_ros_gc
xrc_wwl_7_14 wwl_7_13 wwl_7_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_14 wbl_6_14 wbl_7_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_14 rwl_7_13 rwl_7_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_14 rbl_6_14 rbl_7_14 rc_unit R0=Rrbl C0=Crbl
xgc_7_15 wwl_7_15 wbl_7_15 rwl_7_15 rbl_7_15 sn_7_15 wos_ros_gc
xrc_wwl_7_15 wwl_7_14 wwl_7_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_15 wbl_6_15 wbl_7_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_15 rwl_7_14 rwl_7_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_15 rbl_6_15 rbl_7_15 rc_unit R0=Rrbl C0=Crbl
xgc_7_16 wwl_7_16 wbl_7_16 rwl_7_16 rbl_7_16 sn_7_16 wos_ros_gc
xrc_wwl_7_16 wwl_7_15 wwl_7_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_16 wbl_6_16 wbl_7_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_16 rwl_7_15 rwl_7_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_16 rbl_6_16 rbl_7_16 rc_unit R0=Rrbl C0=Crbl
xgc_7_17 wwl_7_17 wbl_7_17 rwl_7_17 rbl_7_17 sn_7_17 wos_ros_gc
xrc_wwl_7_17 wwl_7_16 wwl_7_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_17 wbl_6_17 wbl_7_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_17 rwl_7_16 rwl_7_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_17 rbl_6_17 rbl_7_17 rc_unit R0=Rrbl C0=Crbl
xgc_7_18 wwl_7_18 wbl_7_18 rwl_7_18 rbl_7_18 sn_7_18 wos_ros_gc
xrc_wwl_7_18 wwl_7_17 wwl_7_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_18 wbl_6_18 wbl_7_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_18 rwl_7_17 rwl_7_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_18 rbl_6_18 rbl_7_18 rc_unit R0=Rrbl C0=Crbl
xgc_7_19 wwl_7_19 wbl_7_19 rwl_7_19 rbl_7_19 sn_7_19 wos_ros_gc
xrc_wwl_7_19 wwl_7_18 wwl_7_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_19 wbl_6_19 wbl_7_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_19 rwl_7_18 rwl_7_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_19 rbl_6_19 rbl_7_19 rc_unit R0=Rrbl C0=Crbl
xgc_7_20 wwl_7_20 wbl_7_20 rwl_7_20 rbl_7_20 sn_7_20 wos_ros_gc
xrc_wwl_7_20 wwl_7_19 wwl_7_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_20 wbl_6_20 wbl_7_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_20 rwl_7_19 rwl_7_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_20 rbl_6_20 rbl_7_20 rc_unit R0=Rrbl C0=Crbl
xgc_7_21 wwl_7_21 wbl_7_21 rwl_7_21 rbl_7_21 sn_7_21 wos_ros_gc
xrc_wwl_7_21 wwl_7_20 wwl_7_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_21 wbl_6_21 wbl_7_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_21 rwl_7_20 rwl_7_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_21 rbl_6_21 rbl_7_21 rc_unit R0=Rrbl C0=Crbl
xgc_7_22 wwl_7_22 wbl_7_22 rwl_7_22 rbl_7_22 sn_7_22 wos_ros_gc
xrc_wwl_7_22 wwl_7_21 wwl_7_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_22 wbl_6_22 wbl_7_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_22 rwl_7_21 rwl_7_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_22 rbl_6_22 rbl_7_22 rc_unit R0=Rrbl C0=Crbl
xgc_7_23 wwl_7_23 wbl_7_23 rwl_7_23 rbl_7_23 sn_7_23 wos_ros_gc
xrc_wwl_7_23 wwl_7_22 wwl_7_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_23 wbl_6_23 wbl_7_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_23 rwl_7_22 rwl_7_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_23 rbl_6_23 rbl_7_23 rc_unit R0=Rrbl C0=Crbl
xgc_7_24 wwl_7_24 wbl_7_24 rwl_7_24 rbl_7_24 sn_7_24 wos_ros_gc
xrc_wwl_7_24 wwl_7_23 wwl_7_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_24 wbl_6_24 wbl_7_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_24 rwl_7_23 rwl_7_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_24 rbl_6_24 rbl_7_24 rc_unit R0=Rrbl C0=Crbl
xgc_7_25 wwl_7_25 wbl_7_25 rwl_7_25 rbl_7_25 sn_7_25 wos_ros_gc
xrc_wwl_7_25 wwl_7_24 wwl_7_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_25 wbl_6_25 wbl_7_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_25 rwl_7_24 rwl_7_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_25 rbl_6_25 rbl_7_25 rc_unit R0=Rrbl C0=Crbl
xgc_7_26 wwl_7_26 wbl_7_26 rwl_7_26 rbl_7_26 sn_7_26 wos_ros_gc
xrc_wwl_7_26 wwl_7_25 wwl_7_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_26 wbl_6_26 wbl_7_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_26 rwl_7_25 rwl_7_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_26 rbl_6_26 rbl_7_26 rc_unit R0=Rrbl C0=Crbl
xgc_7_27 wwl_7_27 wbl_7_27 rwl_7_27 rbl_7_27 sn_7_27 wos_ros_gc
xrc_wwl_7_27 wwl_7_26 wwl_7_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_27 wbl_6_27 wbl_7_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_27 rwl_7_26 rwl_7_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_27 rbl_6_27 rbl_7_27 rc_unit R0=Rrbl C0=Crbl
xgc_7_28 wwl_7_28 wbl_7_28 rwl_7_28 rbl_7_28 sn_7_28 wos_ros_gc
xrc_wwl_7_28 wwl_7_27 wwl_7_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_28 wbl_6_28 wbl_7_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_28 rwl_7_27 rwl_7_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_28 rbl_6_28 rbl_7_28 rc_unit R0=Rrbl C0=Crbl
xgc_7_29 wwl_7_29 wbl_7_29 rwl_7_29 rbl_7_29 sn_7_29 wos_ros_gc
xrc_wwl_7_29 wwl_7_28 wwl_7_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_29 wbl_6_29 wbl_7_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_29 rwl_7_28 rwl_7_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_29 rbl_6_29 rbl_7_29 rc_unit R0=Rrbl C0=Crbl
xgc_7_30 wwl_7_30 wbl_7_30 rwl_7_30 rbl_7_30 sn_7_30 wos_ros_gc
xrc_wwl_7_30 wwl_7_29 wwl_7_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_30 wbl_6_30 wbl_7_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_30 rwl_7_29 rwl_7_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_30 rbl_6_30 rbl_7_30 rc_unit R0=Rrbl C0=Crbl
xgc_7_31 wwl_7_31 wbl_7_31 rwl_7_31 rbl_7_31 sn_7_31 wos_ros_gc
xrc_wwl_7_31 wwl_7_30 wwl_7_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_7_31 wbl_6_31 wbl_7_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_7_31 rwl_7_30 rwl_7_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_7_31 rbl_6_31 rbl_7_31 rc_unit R0=Rrbl C0=Crbl
xgc_8_0 wwl_8_0 wbl_8_0 rwl_8_0 rbl_8_0 sn_8_0 wos_ros_gc
xrc_wwl_8_0 wwl_8 wwl_8_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_0 wbl_7_0 wbl_8_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_0 rwl_8 rwl_8_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_0 rbl_7_0 rbl_8_0 rc_unit R0=Rrbl C0=Crbl
xgc_8_1 wwl_8_1 wbl_8_1 rwl_8_1 rbl_8_1 sn_8_1 wos_ros_gc
xrc_wwl_8_1 wwl_8_0 wwl_8_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_1 wbl_7_1 wbl_8_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_1 rwl_8_0 rwl_8_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_1 rbl_7_1 rbl_8_1 rc_unit R0=Rrbl C0=Crbl
xgc_8_2 wwl_8_2 wbl_8_2 rwl_8_2 rbl_8_2 sn_8_2 wos_ros_gc
xrc_wwl_8_2 wwl_8_1 wwl_8_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_2 wbl_7_2 wbl_8_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_2 rwl_8_1 rwl_8_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_2 rbl_7_2 rbl_8_2 rc_unit R0=Rrbl C0=Crbl
xgc_8_3 wwl_8_3 wbl_8_3 rwl_8_3 rbl_8_3 sn_8_3 wos_ros_gc
xrc_wwl_8_3 wwl_8_2 wwl_8_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_3 wbl_7_3 wbl_8_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_3 rwl_8_2 rwl_8_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_3 rbl_7_3 rbl_8_3 rc_unit R0=Rrbl C0=Crbl
xgc_8_4 wwl_8_4 wbl_8_4 rwl_8_4 rbl_8_4 sn_8_4 wos_ros_gc
xrc_wwl_8_4 wwl_8_3 wwl_8_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_4 wbl_7_4 wbl_8_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_4 rwl_8_3 rwl_8_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_4 rbl_7_4 rbl_8_4 rc_unit R0=Rrbl C0=Crbl
xgc_8_5 wwl_8_5 wbl_8_5 rwl_8_5 rbl_8_5 sn_8_5 wos_ros_gc
xrc_wwl_8_5 wwl_8_4 wwl_8_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_5 wbl_7_5 wbl_8_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_5 rwl_8_4 rwl_8_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_5 rbl_7_5 rbl_8_5 rc_unit R0=Rrbl C0=Crbl
xgc_8_6 wwl_8_6 wbl_8_6 rwl_8_6 rbl_8_6 sn_8_6 wos_ros_gc
xrc_wwl_8_6 wwl_8_5 wwl_8_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_6 wbl_7_6 wbl_8_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_6 rwl_8_5 rwl_8_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_6 rbl_7_6 rbl_8_6 rc_unit R0=Rrbl C0=Crbl
xgc_8_7 wwl_8_7 wbl_8_7 rwl_8_7 rbl_8_7 sn_8_7 wos_ros_gc
xrc_wwl_8_7 wwl_8_6 wwl_8_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_7 wbl_7_7 wbl_8_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_7 rwl_8_6 rwl_8_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_7 rbl_7_7 rbl_8_7 rc_unit R0=Rrbl C0=Crbl
xgc_8_8 wwl_8_8 wbl_8_8 rwl_8_8 rbl_8_8 sn_8_8 wos_ros_gc
xrc_wwl_8_8 wwl_8_7 wwl_8_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_8 wbl_7_8 wbl_8_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_8 rwl_8_7 rwl_8_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_8 rbl_7_8 rbl_8_8 rc_unit R0=Rrbl C0=Crbl
xgc_8_9 wwl_8_9 wbl_8_9 rwl_8_9 rbl_8_9 sn_8_9 wos_ros_gc
xrc_wwl_8_9 wwl_8_8 wwl_8_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_9 wbl_7_9 wbl_8_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_9 rwl_8_8 rwl_8_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_9 rbl_7_9 rbl_8_9 rc_unit R0=Rrbl C0=Crbl
xgc_8_10 wwl_8_10 wbl_8_10 rwl_8_10 rbl_8_10 sn_8_10 wos_ros_gc
xrc_wwl_8_10 wwl_8_9 wwl_8_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_10 wbl_7_10 wbl_8_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_10 rwl_8_9 rwl_8_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_10 rbl_7_10 rbl_8_10 rc_unit R0=Rrbl C0=Crbl
xgc_8_11 wwl_8_11 wbl_8_11 rwl_8_11 rbl_8_11 sn_8_11 wos_ros_gc
xrc_wwl_8_11 wwl_8_10 wwl_8_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_11 wbl_7_11 wbl_8_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_11 rwl_8_10 rwl_8_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_11 rbl_7_11 rbl_8_11 rc_unit R0=Rrbl C0=Crbl
xgc_8_12 wwl_8_12 wbl_8_12 rwl_8_12 rbl_8_12 sn_8_12 wos_ros_gc
xrc_wwl_8_12 wwl_8_11 wwl_8_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_12 wbl_7_12 wbl_8_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_12 rwl_8_11 rwl_8_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_12 rbl_7_12 rbl_8_12 rc_unit R0=Rrbl C0=Crbl
xgc_8_13 wwl_8_13 wbl_8_13 rwl_8_13 rbl_8_13 sn_8_13 wos_ros_gc
xrc_wwl_8_13 wwl_8_12 wwl_8_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_13 wbl_7_13 wbl_8_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_13 rwl_8_12 rwl_8_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_13 rbl_7_13 rbl_8_13 rc_unit R0=Rrbl C0=Crbl
xgc_8_14 wwl_8_14 wbl_8_14 rwl_8_14 rbl_8_14 sn_8_14 wos_ros_gc
xrc_wwl_8_14 wwl_8_13 wwl_8_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_14 wbl_7_14 wbl_8_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_14 rwl_8_13 rwl_8_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_14 rbl_7_14 rbl_8_14 rc_unit R0=Rrbl C0=Crbl
xgc_8_15 wwl_8_15 wbl_8_15 rwl_8_15 rbl_8_15 sn_8_15 wos_ros_gc
xrc_wwl_8_15 wwl_8_14 wwl_8_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_15 wbl_7_15 wbl_8_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_15 rwl_8_14 rwl_8_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_15 rbl_7_15 rbl_8_15 rc_unit R0=Rrbl C0=Crbl
xgc_8_16 wwl_8_16 wbl_8_16 rwl_8_16 rbl_8_16 sn_8_16 wos_ros_gc
xrc_wwl_8_16 wwl_8_15 wwl_8_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_16 wbl_7_16 wbl_8_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_16 rwl_8_15 rwl_8_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_16 rbl_7_16 rbl_8_16 rc_unit R0=Rrbl C0=Crbl
xgc_8_17 wwl_8_17 wbl_8_17 rwl_8_17 rbl_8_17 sn_8_17 wos_ros_gc
xrc_wwl_8_17 wwl_8_16 wwl_8_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_17 wbl_7_17 wbl_8_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_17 rwl_8_16 rwl_8_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_17 rbl_7_17 rbl_8_17 rc_unit R0=Rrbl C0=Crbl
xgc_8_18 wwl_8_18 wbl_8_18 rwl_8_18 rbl_8_18 sn_8_18 wos_ros_gc
xrc_wwl_8_18 wwl_8_17 wwl_8_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_18 wbl_7_18 wbl_8_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_18 rwl_8_17 rwl_8_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_18 rbl_7_18 rbl_8_18 rc_unit R0=Rrbl C0=Crbl
xgc_8_19 wwl_8_19 wbl_8_19 rwl_8_19 rbl_8_19 sn_8_19 wos_ros_gc
xrc_wwl_8_19 wwl_8_18 wwl_8_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_19 wbl_7_19 wbl_8_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_19 rwl_8_18 rwl_8_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_19 rbl_7_19 rbl_8_19 rc_unit R0=Rrbl C0=Crbl
xgc_8_20 wwl_8_20 wbl_8_20 rwl_8_20 rbl_8_20 sn_8_20 wos_ros_gc
xrc_wwl_8_20 wwl_8_19 wwl_8_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_20 wbl_7_20 wbl_8_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_20 rwl_8_19 rwl_8_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_20 rbl_7_20 rbl_8_20 rc_unit R0=Rrbl C0=Crbl
xgc_8_21 wwl_8_21 wbl_8_21 rwl_8_21 rbl_8_21 sn_8_21 wos_ros_gc
xrc_wwl_8_21 wwl_8_20 wwl_8_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_21 wbl_7_21 wbl_8_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_21 rwl_8_20 rwl_8_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_21 rbl_7_21 rbl_8_21 rc_unit R0=Rrbl C0=Crbl
xgc_8_22 wwl_8_22 wbl_8_22 rwl_8_22 rbl_8_22 sn_8_22 wos_ros_gc
xrc_wwl_8_22 wwl_8_21 wwl_8_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_22 wbl_7_22 wbl_8_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_22 rwl_8_21 rwl_8_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_22 rbl_7_22 rbl_8_22 rc_unit R0=Rrbl C0=Crbl
xgc_8_23 wwl_8_23 wbl_8_23 rwl_8_23 rbl_8_23 sn_8_23 wos_ros_gc
xrc_wwl_8_23 wwl_8_22 wwl_8_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_23 wbl_7_23 wbl_8_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_23 rwl_8_22 rwl_8_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_23 rbl_7_23 rbl_8_23 rc_unit R0=Rrbl C0=Crbl
xgc_8_24 wwl_8_24 wbl_8_24 rwl_8_24 rbl_8_24 sn_8_24 wos_ros_gc
xrc_wwl_8_24 wwl_8_23 wwl_8_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_24 wbl_7_24 wbl_8_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_24 rwl_8_23 rwl_8_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_24 rbl_7_24 rbl_8_24 rc_unit R0=Rrbl C0=Crbl
xgc_8_25 wwl_8_25 wbl_8_25 rwl_8_25 rbl_8_25 sn_8_25 wos_ros_gc
xrc_wwl_8_25 wwl_8_24 wwl_8_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_25 wbl_7_25 wbl_8_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_25 rwl_8_24 rwl_8_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_25 rbl_7_25 rbl_8_25 rc_unit R0=Rrbl C0=Crbl
xgc_8_26 wwl_8_26 wbl_8_26 rwl_8_26 rbl_8_26 sn_8_26 wos_ros_gc
xrc_wwl_8_26 wwl_8_25 wwl_8_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_26 wbl_7_26 wbl_8_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_26 rwl_8_25 rwl_8_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_26 rbl_7_26 rbl_8_26 rc_unit R0=Rrbl C0=Crbl
xgc_8_27 wwl_8_27 wbl_8_27 rwl_8_27 rbl_8_27 sn_8_27 wos_ros_gc
xrc_wwl_8_27 wwl_8_26 wwl_8_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_27 wbl_7_27 wbl_8_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_27 rwl_8_26 rwl_8_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_27 rbl_7_27 rbl_8_27 rc_unit R0=Rrbl C0=Crbl
xgc_8_28 wwl_8_28 wbl_8_28 rwl_8_28 rbl_8_28 sn_8_28 wos_ros_gc
xrc_wwl_8_28 wwl_8_27 wwl_8_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_28 wbl_7_28 wbl_8_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_28 rwl_8_27 rwl_8_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_28 rbl_7_28 rbl_8_28 rc_unit R0=Rrbl C0=Crbl
xgc_8_29 wwl_8_29 wbl_8_29 rwl_8_29 rbl_8_29 sn_8_29 wos_ros_gc
xrc_wwl_8_29 wwl_8_28 wwl_8_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_29 wbl_7_29 wbl_8_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_29 rwl_8_28 rwl_8_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_29 rbl_7_29 rbl_8_29 rc_unit R0=Rrbl C0=Crbl
xgc_8_30 wwl_8_30 wbl_8_30 rwl_8_30 rbl_8_30 sn_8_30 wos_ros_gc
xrc_wwl_8_30 wwl_8_29 wwl_8_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_30 wbl_7_30 wbl_8_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_30 rwl_8_29 rwl_8_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_30 rbl_7_30 rbl_8_30 rc_unit R0=Rrbl C0=Crbl
xgc_8_31 wwl_8_31 wbl_8_31 rwl_8_31 rbl_8_31 sn_8_31 wos_ros_gc
xrc_wwl_8_31 wwl_8_30 wwl_8_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_8_31 wbl_7_31 wbl_8_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_8_31 rwl_8_30 rwl_8_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_8_31 rbl_7_31 rbl_8_31 rc_unit R0=Rrbl C0=Crbl
xgc_9_0 wwl_9_0 wbl_9_0 rwl_9_0 rbl_9_0 sn_9_0 wos_ros_gc
xrc_wwl_9_0 wwl_9 wwl_9_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_0 wbl_8_0 wbl_9_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_0 rwl_9 rwl_9_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_0 rbl_8_0 rbl_9_0 rc_unit R0=Rrbl C0=Crbl
xgc_9_1 wwl_9_1 wbl_9_1 rwl_9_1 rbl_9_1 sn_9_1 wos_ros_gc
xrc_wwl_9_1 wwl_9_0 wwl_9_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_1 wbl_8_1 wbl_9_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_1 rwl_9_0 rwl_9_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_1 rbl_8_1 rbl_9_1 rc_unit R0=Rrbl C0=Crbl
xgc_9_2 wwl_9_2 wbl_9_2 rwl_9_2 rbl_9_2 sn_9_2 wos_ros_gc
xrc_wwl_9_2 wwl_9_1 wwl_9_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_2 wbl_8_2 wbl_9_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_2 rwl_9_1 rwl_9_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_2 rbl_8_2 rbl_9_2 rc_unit R0=Rrbl C0=Crbl
xgc_9_3 wwl_9_3 wbl_9_3 rwl_9_3 rbl_9_3 sn_9_3 wos_ros_gc
xrc_wwl_9_3 wwl_9_2 wwl_9_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_3 wbl_8_3 wbl_9_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_3 rwl_9_2 rwl_9_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_3 rbl_8_3 rbl_9_3 rc_unit R0=Rrbl C0=Crbl
xgc_9_4 wwl_9_4 wbl_9_4 rwl_9_4 rbl_9_4 sn_9_4 wos_ros_gc
xrc_wwl_9_4 wwl_9_3 wwl_9_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_4 wbl_8_4 wbl_9_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_4 rwl_9_3 rwl_9_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_4 rbl_8_4 rbl_9_4 rc_unit R0=Rrbl C0=Crbl
xgc_9_5 wwl_9_5 wbl_9_5 rwl_9_5 rbl_9_5 sn_9_5 wos_ros_gc
xrc_wwl_9_5 wwl_9_4 wwl_9_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_5 wbl_8_5 wbl_9_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_5 rwl_9_4 rwl_9_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_5 rbl_8_5 rbl_9_5 rc_unit R0=Rrbl C0=Crbl
xgc_9_6 wwl_9_6 wbl_9_6 rwl_9_6 rbl_9_6 sn_9_6 wos_ros_gc
xrc_wwl_9_6 wwl_9_5 wwl_9_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_6 wbl_8_6 wbl_9_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_6 rwl_9_5 rwl_9_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_6 rbl_8_6 rbl_9_6 rc_unit R0=Rrbl C0=Crbl
xgc_9_7 wwl_9_7 wbl_9_7 rwl_9_7 rbl_9_7 sn_9_7 wos_ros_gc
xrc_wwl_9_7 wwl_9_6 wwl_9_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_7 wbl_8_7 wbl_9_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_7 rwl_9_6 rwl_9_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_7 rbl_8_7 rbl_9_7 rc_unit R0=Rrbl C0=Crbl
xgc_9_8 wwl_9_8 wbl_9_8 rwl_9_8 rbl_9_8 sn_9_8 wos_ros_gc
xrc_wwl_9_8 wwl_9_7 wwl_9_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_8 wbl_8_8 wbl_9_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_8 rwl_9_7 rwl_9_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_8 rbl_8_8 rbl_9_8 rc_unit R0=Rrbl C0=Crbl
xgc_9_9 wwl_9_9 wbl_9_9 rwl_9_9 rbl_9_9 sn_9_9 wos_ros_gc
xrc_wwl_9_9 wwl_9_8 wwl_9_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_9 wbl_8_9 wbl_9_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_9 rwl_9_8 rwl_9_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_9 rbl_8_9 rbl_9_9 rc_unit R0=Rrbl C0=Crbl
xgc_9_10 wwl_9_10 wbl_9_10 rwl_9_10 rbl_9_10 sn_9_10 wos_ros_gc
xrc_wwl_9_10 wwl_9_9 wwl_9_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_10 wbl_8_10 wbl_9_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_10 rwl_9_9 rwl_9_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_10 rbl_8_10 rbl_9_10 rc_unit R0=Rrbl C0=Crbl
xgc_9_11 wwl_9_11 wbl_9_11 rwl_9_11 rbl_9_11 sn_9_11 wos_ros_gc
xrc_wwl_9_11 wwl_9_10 wwl_9_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_11 wbl_8_11 wbl_9_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_11 rwl_9_10 rwl_9_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_11 rbl_8_11 rbl_9_11 rc_unit R0=Rrbl C0=Crbl
xgc_9_12 wwl_9_12 wbl_9_12 rwl_9_12 rbl_9_12 sn_9_12 wos_ros_gc
xrc_wwl_9_12 wwl_9_11 wwl_9_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_12 wbl_8_12 wbl_9_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_12 rwl_9_11 rwl_9_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_12 rbl_8_12 rbl_9_12 rc_unit R0=Rrbl C0=Crbl
xgc_9_13 wwl_9_13 wbl_9_13 rwl_9_13 rbl_9_13 sn_9_13 wos_ros_gc
xrc_wwl_9_13 wwl_9_12 wwl_9_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_13 wbl_8_13 wbl_9_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_13 rwl_9_12 rwl_9_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_13 rbl_8_13 rbl_9_13 rc_unit R0=Rrbl C0=Crbl
xgc_9_14 wwl_9_14 wbl_9_14 rwl_9_14 rbl_9_14 sn_9_14 wos_ros_gc
xrc_wwl_9_14 wwl_9_13 wwl_9_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_14 wbl_8_14 wbl_9_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_14 rwl_9_13 rwl_9_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_14 rbl_8_14 rbl_9_14 rc_unit R0=Rrbl C0=Crbl
xgc_9_15 wwl_9_15 wbl_9_15 rwl_9_15 rbl_9_15 sn_9_15 wos_ros_gc
xrc_wwl_9_15 wwl_9_14 wwl_9_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_15 wbl_8_15 wbl_9_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_15 rwl_9_14 rwl_9_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_15 rbl_8_15 rbl_9_15 rc_unit R0=Rrbl C0=Crbl
xgc_9_16 wwl_9_16 wbl_9_16 rwl_9_16 rbl_9_16 sn_9_16 wos_ros_gc
xrc_wwl_9_16 wwl_9_15 wwl_9_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_16 wbl_8_16 wbl_9_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_16 rwl_9_15 rwl_9_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_16 rbl_8_16 rbl_9_16 rc_unit R0=Rrbl C0=Crbl
xgc_9_17 wwl_9_17 wbl_9_17 rwl_9_17 rbl_9_17 sn_9_17 wos_ros_gc
xrc_wwl_9_17 wwl_9_16 wwl_9_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_17 wbl_8_17 wbl_9_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_17 rwl_9_16 rwl_9_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_17 rbl_8_17 rbl_9_17 rc_unit R0=Rrbl C0=Crbl
xgc_9_18 wwl_9_18 wbl_9_18 rwl_9_18 rbl_9_18 sn_9_18 wos_ros_gc
xrc_wwl_9_18 wwl_9_17 wwl_9_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_18 wbl_8_18 wbl_9_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_18 rwl_9_17 rwl_9_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_18 rbl_8_18 rbl_9_18 rc_unit R0=Rrbl C0=Crbl
xgc_9_19 wwl_9_19 wbl_9_19 rwl_9_19 rbl_9_19 sn_9_19 wos_ros_gc
xrc_wwl_9_19 wwl_9_18 wwl_9_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_19 wbl_8_19 wbl_9_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_19 rwl_9_18 rwl_9_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_19 rbl_8_19 rbl_9_19 rc_unit R0=Rrbl C0=Crbl
xgc_9_20 wwl_9_20 wbl_9_20 rwl_9_20 rbl_9_20 sn_9_20 wos_ros_gc
xrc_wwl_9_20 wwl_9_19 wwl_9_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_20 wbl_8_20 wbl_9_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_20 rwl_9_19 rwl_9_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_20 rbl_8_20 rbl_9_20 rc_unit R0=Rrbl C0=Crbl
xgc_9_21 wwl_9_21 wbl_9_21 rwl_9_21 rbl_9_21 sn_9_21 wos_ros_gc
xrc_wwl_9_21 wwl_9_20 wwl_9_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_21 wbl_8_21 wbl_9_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_21 rwl_9_20 rwl_9_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_21 rbl_8_21 rbl_9_21 rc_unit R0=Rrbl C0=Crbl
xgc_9_22 wwl_9_22 wbl_9_22 rwl_9_22 rbl_9_22 sn_9_22 wos_ros_gc
xrc_wwl_9_22 wwl_9_21 wwl_9_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_22 wbl_8_22 wbl_9_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_22 rwl_9_21 rwl_9_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_22 rbl_8_22 rbl_9_22 rc_unit R0=Rrbl C0=Crbl
xgc_9_23 wwl_9_23 wbl_9_23 rwl_9_23 rbl_9_23 sn_9_23 wos_ros_gc
xrc_wwl_9_23 wwl_9_22 wwl_9_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_23 wbl_8_23 wbl_9_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_23 rwl_9_22 rwl_9_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_23 rbl_8_23 rbl_9_23 rc_unit R0=Rrbl C0=Crbl
xgc_9_24 wwl_9_24 wbl_9_24 rwl_9_24 rbl_9_24 sn_9_24 wos_ros_gc
xrc_wwl_9_24 wwl_9_23 wwl_9_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_24 wbl_8_24 wbl_9_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_24 rwl_9_23 rwl_9_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_24 rbl_8_24 rbl_9_24 rc_unit R0=Rrbl C0=Crbl
xgc_9_25 wwl_9_25 wbl_9_25 rwl_9_25 rbl_9_25 sn_9_25 wos_ros_gc
xrc_wwl_9_25 wwl_9_24 wwl_9_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_25 wbl_8_25 wbl_9_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_25 rwl_9_24 rwl_9_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_25 rbl_8_25 rbl_9_25 rc_unit R0=Rrbl C0=Crbl
xgc_9_26 wwl_9_26 wbl_9_26 rwl_9_26 rbl_9_26 sn_9_26 wos_ros_gc
xrc_wwl_9_26 wwl_9_25 wwl_9_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_26 wbl_8_26 wbl_9_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_26 rwl_9_25 rwl_9_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_26 rbl_8_26 rbl_9_26 rc_unit R0=Rrbl C0=Crbl
xgc_9_27 wwl_9_27 wbl_9_27 rwl_9_27 rbl_9_27 sn_9_27 wos_ros_gc
xrc_wwl_9_27 wwl_9_26 wwl_9_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_27 wbl_8_27 wbl_9_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_27 rwl_9_26 rwl_9_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_27 rbl_8_27 rbl_9_27 rc_unit R0=Rrbl C0=Crbl
xgc_9_28 wwl_9_28 wbl_9_28 rwl_9_28 rbl_9_28 sn_9_28 wos_ros_gc
xrc_wwl_9_28 wwl_9_27 wwl_9_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_28 wbl_8_28 wbl_9_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_28 rwl_9_27 rwl_9_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_28 rbl_8_28 rbl_9_28 rc_unit R0=Rrbl C0=Crbl
xgc_9_29 wwl_9_29 wbl_9_29 rwl_9_29 rbl_9_29 sn_9_29 wos_ros_gc
xrc_wwl_9_29 wwl_9_28 wwl_9_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_29 wbl_8_29 wbl_9_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_29 rwl_9_28 rwl_9_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_29 rbl_8_29 rbl_9_29 rc_unit R0=Rrbl C0=Crbl
xgc_9_30 wwl_9_30 wbl_9_30 rwl_9_30 rbl_9_30 sn_9_30 wos_ros_gc
xrc_wwl_9_30 wwl_9_29 wwl_9_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_30 wbl_8_30 wbl_9_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_30 rwl_9_29 rwl_9_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_30 rbl_8_30 rbl_9_30 rc_unit R0=Rrbl C0=Crbl
xgc_9_31 wwl_9_31 wbl_9_31 rwl_9_31 rbl_9_31 sn_9_31 wos_ros_gc
xrc_wwl_9_31 wwl_9_30 wwl_9_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_9_31 wbl_8_31 wbl_9_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_9_31 rwl_9_30 rwl_9_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_9_31 rbl_8_31 rbl_9_31 rc_unit R0=Rrbl C0=Crbl
xgc_10_0 wwl_10_0 wbl_10_0 rwl_10_0 rbl_10_0 sn_10_0 wos_ros_gc
xrc_wwl_10_0 wwl_10 wwl_10_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_0 wbl_9_0 wbl_10_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_0 rwl_10 rwl_10_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_0 rbl_9_0 rbl_10_0 rc_unit R0=Rrbl C0=Crbl
xgc_10_1 wwl_10_1 wbl_10_1 rwl_10_1 rbl_10_1 sn_10_1 wos_ros_gc
xrc_wwl_10_1 wwl_10_0 wwl_10_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_1 wbl_9_1 wbl_10_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_1 rwl_10_0 rwl_10_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_1 rbl_9_1 rbl_10_1 rc_unit R0=Rrbl C0=Crbl
xgc_10_2 wwl_10_2 wbl_10_2 rwl_10_2 rbl_10_2 sn_10_2 wos_ros_gc
xrc_wwl_10_2 wwl_10_1 wwl_10_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_2 wbl_9_2 wbl_10_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_2 rwl_10_1 rwl_10_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_2 rbl_9_2 rbl_10_2 rc_unit R0=Rrbl C0=Crbl
xgc_10_3 wwl_10_3 wbl_10_3 rwl_10_3 rbl_10_3 sn_10_3 wos_ros_gc
xrc_wwl_10_3 wwl_10_2 wwl_10_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_3 wbl_9_3 wbl_10_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_3 rwl_10_2 rwl_10_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_3 rbl_9_3 rbl_10_3 rc_unit R0=Rrbl C0=Crbl
xgc_10_4 wwl_10_4 wbl_10_4 rwl_10_4 rbl_10_4 sn_10_4 wos_ros_gc
xrc_wwl_10_4 wwl_10_3 wwl_10_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_4 wbl_9_4 wbl_10_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_4 rwl_10_3 rwl_10_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_4 rbl_9_4 rbl_10_4 rc_unit R0=Rrbl C0=Crbl
xgc_10_5 wwl_10_5 wbl_10_5 rwl_10_5 rbl_10_5 sn_10_5 wos_ros_gc
xrc_wwl_10_5 wwl_10_4 wwl_10_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_5 wbl_9_5 wbl_10_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_5 rwl_10_4 rwl_10_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_5 rbl_9_5 rbl_10_5 rc_unit R0=Rrbl C0=Crbl
xgc_10_6 wwl_10_6 wbl_10_6 rwl_10_6 rbl_10_6 sn_10_6 wos_ros_gc
xrc_wwl_10_6 wwl_10_5 wwl_10_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_6 wbl_9_6 wbl_10_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_6 rwl_10_5 rwl_10_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_6 rbl_9_6 rbl_10_6 rc_unit R0=Rrbl C0=Crbl
xgc_10_7 wwl_10_7 wbl_10_7 rwl_10_7 rbl_10_7 sn_10_7 wos_ros_gc
xrc_wwl_10_7 wwl_10_6 wwl_10_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_7 wbl_9_7 wbl_10_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_7 rwl_10_6 rwl_10_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_7 rbl_9_7 rbl_10_7 rc_unit R0=Rrbl C0=Crbl
xgc_10_8 wwl_10_8 wbl_10_8 rwl_10_8 rbl_10_8 sn_10_8 wos_ros_gc
xrc_wwl_10_8 wwl_10_7 wwl_10_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_8 wbl_9_8 wbl_10_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_8 rwl_10_7 rwl_10_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_8 rbl_9_8 rbl_10_8 rc_unit R0=Rrbl C0=Crbl
xgc_10_9 wwl_10_9 wbl_10_9 rwl_10_9 rbl_10_9 sn_10_9 wos_ros_gc
xrc_wwl_10_9 wwl_10_8 wwl_10_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_9 wbl_9_9 wbl_10_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_9 rwl_10_8 rwl_10_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_9 rbl_9_9 rbl_10_9 rc_unit R0=Rrbl C0=Crbl
xgc_10_10 wwl_10_10 wbl_10_10 rwl_10_10 rbl_10_10 sn_10_10 wos_ros_gc
xrc_wwl_10_10 wwl_10_9 wwl_10_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_10 wbl_9_10 wbl_10_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_10 rwl_10_9 rwl_10_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_10 rbl_9_10 rbl_10_10 rc_unit R0=Rrbl C0=Crbl
xgc_10_11 wwl_10_11 wbl_10_11 rwl_10_11 rbl_10_11 sn_10_11 wos_ros_gc
xrc_wwl_10_11 wwl_10_10 wwl_10_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_11 wbl_9_11 wbl_10_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_11 rwl_10_10 rwl_10_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_11 rbl_9_11 rbl_10_11 rc_unit R0=Rrbl C0=Crbl
xgc_10_12 wwl_10_12 wbl_10_12 rwl_10_12 rbl_10_12 sn_10_12 wos_ros_gc
xrc_wwl_10_12 wwl_10_11 wwl_10_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_12 wbl_9_12 wbl_10_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_12 rwl_10_11 rwl_10_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_12 rbl_9_12 rbl_10_12 rc_unit R0=Rrbl C0=Crbl
xgc_10_13 wwl_10_13 wbl_10_13 rwl_10_13 rbl_10_13 sn_10_13 wos_ros_gc
xrc_wwl_10_13 wwl_10_12 wwl_10_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_13 wbl_9_13 wbl_10_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_13 rwl_10_12 rwl_10_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_13 rbl_9_13 rbl_10_13 rc_unit R0=Rrbl C0=Crbl
xgc_10_14 wwl_10_14 wbl_10_14 rwl_10_14 rbl_10_14 sn_10_14 wos_ros_gc
xrc_wwl_10_14 wwl_10_13 wwl_10_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_14 wbl_9_14 wbl_10_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_14 rwl_10_13 rwl_10_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_14 rbl_9_14 rbl_10_14 rc_unit R0=Rrbl C0=Crbl
xgc_10_15 wwl_10_15 wbl_10_15 rwl_10_15 rbl_10_15 sn_10_15 wos_ros_gc
xrc_wwl_10_15 wwl_10_14 wwl_10_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_15 wbl_9_15 wbl_10_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_15 rwl_10_14 rwl_10_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_15 rbl_9_15 rbl_10_15 rc_unit R0=Rrbl C0=Crbl
xgc_10_16 wwl_10_16 wbl_10_16 rwl_10_16 rbl_10_16 sn_10_16 wos_ros_gc
xrc_wwl_10_16 wwl_10_15 wwl_10_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_16 wbl_9_16 wbl_10_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_16 rwl_10_15 rwl_10_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_16 rbl_9_16 rbl_10_16 rc_unit R0=Rrbl C0=Crbl
xgc_10_17 wwl_10_17 wbl_10_17 rwl_10_17 rbl_10_17 sn_10_17 wos_ros_gc
xrc_wwl_10_17 wwl_10_16 wwl_10_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_17 wbl_9_17 wbl_10_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_17 rwl_10_16 rwl_10_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_17 rbl_9_17 rbl_10_17 rc_unit R0=Rrbl C0=Crbl
xgc_10_18 wwl_10_18 wbl_10_18 rwl_10_18 rbl_10_18 sn_10_18 wos_ros_gc
xrc_wwl_10_18 wwl_10_17 wwl_10_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_18 wbl_9_18 wbl_10_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_18 rwl_10_17 rwl_10_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_18 rbl_9_18 rbl_10_18 rc_unit R0=Rrbl C0=Crbl
xgc_10_19 wwl_10_19 wbl_10_19 rwl_10_19 rbl_10_19 sn_10_19 wos_ros_gc
xrc_wwl_10_19 wwl_10_18 wwl_10_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_19 wbl_9_19 wbl_10_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_19 rwl_10_18 rwl_10_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_19 rbl_9_19 rbl_10_19 rc_unit R0=Rrbl C0=Crbl
xgc_10_20 wwl_10_20 wbl_10_20 rwl_10_20 rbl_10_20 sn_10_20 wos_ros_gc
xrc_wwl_10_20 wwl_10_19 wwl_10_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_20 wbl_9_20 wbl_10_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_20 rwl_10_19 rwl_10_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_20 rbl_9_20 rbl_10_20 rc_unit R0=Rrbl C0=Crbl
xgc_10_21 wwl_10_21 wbl_10_21 rwl_10_21 rbl_10_21 sn_10_21 wos_ros_gc
xrc_wwl_10_21 wwl_10_20 wwl_10_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_21 wbl_9_21 wbl_10_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_21 rwl_10_20 rwl_10_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_21 rbl_9_21 rbl_10_21 rc_unit R0=Rrbl C0=Crbl
xgc_10_22 wwl_10_22 wbl_10_22 rwl_10_22 rbl_10_22 sn_10_22 wos_ros_gc
xrc_wwl_10_22 wwl_10_21 wwl_10_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_22 wbl_9_22 wbl_10_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_22 rwl_10_21 rwl_10_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_22 rbl_9_22 rbl_10_22 rc_unit R0=Rrbl C0=Crbl
xgc_10_23 wwl_10_23 wbl_10_23 rwl_10_23 rbl_10_23 sn_10_23 wos_ros_gc
xrc_wwl_10_23 wwl_10_22 wwl_10_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_23 wbl_9_23 wbl_10_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_23 rwl_10_22 rwl_10_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_23 rbl_9_23 rbl_10_23 rc_unit R0=Rrbl C0=Crbl
xgc_10_24 wwl_10_24 wbl_10_24 rwl_10_24 rbl_10_24 sn_10_24 wos_ros_gc
xrc_wwl_10_24 wwl_10_23 wwl_10_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_24 wbl_9_24 wbl_10_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_24 rwl_10_23 rwl_10_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_24 rbl_9_24 rbl_10_24 rc_unit R0=Rrbl C0=Crbl
xgc_10_25 wwl_10_25 wbl_10_25 rwl_10_25 rbl_10_25 sn_10_25 wos_ros_gc
xrc_wwl_10_25 wwl_10_24 wwl_10_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_25 wbl_9_25 wbl_10_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_25 rwl_10_24 rwl_10_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_25 rbl_9_25 rbl_10_25 rc_unit R0=Rrbl C0=Crbl
xgc_10_26 wwl_10_26 wbl_10_26 rwl_10_26 rbl_10_26 sn_10_26 wos_ros_gc
xrc_wwl_10_26 wwl_10_25 wwl_10_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_26 wbl_9_26 wbl_10_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_26 rwl_10_25 rwl_10_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_26 rbl_9_26 rbl_10_26 rc_unit R0=Rrbl C0=Crbl
xgc_10_27 wwl_10_27 wbl_10_27 rwl_10_27 rbl_10_27 sn_10_27 wos_ros_gc
xrc_wwl_10_27 wwl_10_26 wwl_10_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_27 wbl_9_27 wbl_10_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_27 rwl_10_26 rwl_10_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_27 rbl_9_27 rbl_10_27 rc_unit R0=Rrbl C0=Crbl
xgc_10_28 wwl_10_28 wbl_10_28 rwl_10_28 rbl_10_28 sn_10_28 wos_ros_gc
xrc_wwl_10_28 wwl_10_27 wwl_10_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_28 wbl_9_28 wbl_10_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_28 rwl_10_27 rwl_10_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_28 rbl_9_28 rbl_10_28 rc_unit R0=Rrbl C0=Crbl
xgc_10_29 wwl_10_29 wbl_10_29 rwl_10_29 rbl_10_29 sn_10_29 wos_ros_gc
xrc_wwl_10_29 wwl_10_28 wwl_10_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_29 wbl_9_29 wbl_10_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_29 rwl_10_28 rwl_10_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_29 rbl_9_29 rbl_10_29 rc_unit R0=Rrbl C0=Crbl
xgc_10_30 wwl_10_30 wbl_10_30 rwl_10_30 rbl_10_30 sn_10_30 wos_ros_gc
xrc_wwl_10_30 wwl_10_29 wwl_10_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_30 wbl_9_30 wbl_10_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_30 rwl_10_29 rwl_10_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_30 rbl_9_30 rbl_10_30 rc_unit R0=Rrbl C0=Crbl
xgc_10_31 wwl_10_31 wbl_10_31 rwl_10_31 rbl_10_31 sn_10_31 wos_ros_gc
xrc_wwl_10_31 wwl_10_30 wwl_10_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_10_31 wbl_9_31 wbl_10_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_10_31 rwl_10_30 rwl_10_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_10_31 rbl_9_31 rbl_10_31 rc_unit R0=Rrbl C0=Crbl
xgc_11_0 wwl_11_0 wbl_11_0 rwl_11_0 rbl_11_0 sn_11_0 wos_ros_gc
xrc_wwl_11_0 wwl_11 wwl_11_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_0 wbl_10_0 wbl_11_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_0 rwl_11 rwl_11_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_0 rbl_10_0 rbl_11_0 rc_unit R0=Rrbl C0=Crbl
xgc_11_1 wwl_11_1 wbl_11_1 rwl_11_1 rbl_11_1 sn_11_1 wos_ros_gc
xrc_wwl_11_1 wwl_11_0 wwl_11_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_1 wbl_10_1 wbl_11_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_1 rwl_11_0 rwl_11_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_1 rbl_10_1 rbl_11_1 rc_unit R0=Rrbl C0=Crbl
xgc_11_2 wwl_11_2 wbl_11_2 rwl_11_2 rbl_11_2 sn_11_2 wos_ros_gc
xrc_wwl_11_2 wwl_11_1 wwl_11_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_2 wbl_10_2 wbl_11_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_2 rwl_11_1 rwl_11_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_2 rbl_10_2 rbl_11_2 rc_unit R0=Rrbl C0=Crbl
xgc_11_3 wwl_11_3 wbl_11_3 rwl_11_3 rbl_11_3 sn_11_3 wos_ros_gc
xrc_wwl_11_3 wwl_11_2 wwl_11_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_3 wbl_10_3 wbl_11_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_3 rwl_11_2 rwl_11_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_3 rbl_10_3 rbl_11_3 rc_unit R0=Rrbl C0=Crbl
xgc_11_4 wwl_11_4 wbl_11_4 rwl_11_4 rbl_11_4 sn_11_4 wos_ros_gc
xrc_wwl_11_4 wwl_11_3 wwl_11_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_4 wbl_10_4 wbl_11_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_4 rwl_11_3 rwl_11_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_4 rbl_10_4 rbl_11_4 rc_unit R0=Rrbl C0=Crbl
xgc_11_5 wwl_11_5 wbl_11_5 rwl_11_5 rbl_11_5 sn_11_5 wos_ros_gc
xrc_wwl_11_5 wwl_11_4 wwl_11_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_5 wbl_10_5 wbl_11_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_5 rwl_11_4 rwl_11_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_5 rbl_10_5 rbl_11_5 rc_unit R0=Rrbl C0=Crbl
xgc_11_6 wwl_11_6 wbl_11_6 rwl_11_6 rbl_11_6 sn_11_6 wos_ros_gc
xrc_wwl_11_6 wwl_11_5 wwl_11_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_6 wbl_10_6 wbl_11_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_6 rwl_11_5 rwl_11_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_6 rbl_10_6 rbl_11_6 rc_unit R0=Rrbl C0=Crbl
xgc_11_7 wwl_11_7 wbl_11_7 rwl_11_7 rbl_11_7 sn_11_7 wos_ros_gc
xrc_wwl_11_7 wwl_11_6 wwl_11_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_7 wbl_10_7 wbl_11_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_7 rwl_11_6 rwl_11_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_7 rbl_10_7 rbl_11_7 rc_unit R0=Rrbl C0=Crbl
xgc_11_8 wwl_11_8 wbl_11_8 rwl_11_8 rbl_11_8 sn_11_8 wos_ros_gc
xrc_wwl_11_8 wwl_11_7 wwl_11_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_8 wbl_10_8 wbl_11_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_8 rwl_11_7 rwl_11_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_8 rbl_10_8 rbl_11_8 rc_unit R0=Rrbl C0=Crbl
xgc_11_9 wwl_11_9 wbl_11_9 rwl_11_9 rbl_11_9 sn_11_9 wos_ros_gc
xrc_wwl_11_9 wwl_11_8 wwl_11_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_9 wbl_10_9 wbl_11_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_9 rwl_11_8 rwl_11_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_9 rbl_10_9 rbl_11_9 rc_unit R0=Rrbl C0=Crbl
xgc_11_10 wwl_11_10 wbl_11_10 rwl_11_10 rbl_11_10 sn_11_10 wos_ros_gc
xrc_wwl_11_10 wwl_11_9 wwl_11_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_10 wbl_10_10 wbl_11_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_10 rwl_11_9 rwl_11_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_10 rbl_10_10 rbl_11_10 rc_unit R0=Rrbl C0=Crbl
xgc_11_11 wwl_11_11 wbl_11_11 rwl_11_11 rbl_11_11 sn_11_11 wos_ros_gc
xrc_wwl_11_11 wwl_11_10 wwl_11_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_11 wbl_10_11 wbl_11_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_11 rwl_11_10 rwl_11_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_11 rbl_10_11 rbl_11_11 rc_unit R0=Rrbl C0=Crbl
xgc_11_12 wwl_11_12 wbl_11_12 rwl_11_12 rbl_11_12 sn_11_12 wos_ros_gc
xrc_wwl_11_12 wwl_11_11 wwl_11_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_12 wbl_10_12 wbl_11_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_12 rwl_11_11 rwl_11_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_12 rbl_10_12 rbl_11_12 rc_unit R0=Rrbl C0=Crbl
xgc_11_13 wwl_11_13 wbl_11_13 rwl_11_13 rbl_11_13 sn_11_13 wos_ros_gc
xrc_wwl_11_13 wwl_11_12 wwl_11_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_13 wbl_10_13 wbl_11_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_13 rwl_11_12 rwl_11_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_13 rbl_10_13 rbl_11_13 rc_unit R0=Rrbl C0=Crbl
xgc_11_14 wwl_11_14 wbl_11_14 rwl_11_14 rbl_11_14 sn_11_14 wos_ros_gc
xrc_wwl_11_14 wwl_11_13 wwl_11_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_14 wbl_10_14 wbl_11_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_14 rwl_11_13 rwl_11_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_14 rbl_10_14 rbl_11_14 rc_unit R0=Rrbl C0=Crbl
xgc_11_15 wwl_11_15 wbl_11_15 rwl_11_15 rbl_11_15 sn_11_15 wos_ros_gc
xrc_wwl_11_15 wwl_11_14 wwl_11_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_15 wbl_10_15 wbl_11_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_15 rwl_11_14 rwl_11_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_15 rbl_10_15 rbl_11_15 rc_unit R0=Rrbl C0=Crbl
xgc_11_16 wwl_11_16 wbl_11_16 rwl_11_16 rbl_11_16 sn_11_16 wos_ros_gc
xrc_wwl_11_16 wwl_11_15 wwl_11_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_16 wbl_10_16 wbl_11_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_16 rwl_11_15 rwl_11_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_16 rbl_10_16 rbl_11_16 rc_unit R0=Rrbl C0=Crbl
xgc_11_17 wwl_11_17 wbl_11_17 rwl_11_17 rbl_11_17 sn_11_17 wos_ros_gc
xrc_wwl_11_17 wwl_11_16 wwl_11_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_17 wbl_10_17 wbl_11_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_17 rwl_11_16 rwl_11_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_17 rbl_10_17 rbl_11_17 rc_unit R0=Rrbl C0=Crbl
xgc_11_18 wwl_11_18 wbl_11_18 rwl_11_18 rbl_11_18 sn_11_18 wos_ros_gc
xrc_wwl_11_18 wwl_11_17 wwl_11_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_18 wbl_10_18 wbl_11_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_18 rwl_11_17 rwl_11_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_18 rbl_10_18 rbl_11_18 rc_unit R0=Rrbl C0=Crbl
xgc_11_19 wwl_11_19 wbl_11_19 rwl_11_19 rbl_11_19 sn_11_19 wos_ros_gc
xrc_wwl_11_19 wwl_11_18 wwl_11_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_19 wbl_10_19 wbl_11_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_19 rwl_11_18 rwl_11_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_19 rbl_10_19 rbl_11_19 rc_unit R0=Rrbl C0=Crbl
xgc_11_20 wwl_11_20 wbl_11_20 rwl_11_20 rbl_11_20 sn_11_20 wos_ros_gc
xrc_wwl_11_20 wwl_11_19 wwl_11_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_20 wbl_10_20 wbl_11_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_20 rwl_11_19 rwl_11_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_20 rbl_10_20 rbl_11_20 rc_unit R0=Rrbl C0=Crbl
xgc_11_21 wwl_11_21 wbl_11_21 rwl_11_21 rbl_11_21 sn_11_21 wos_ros_gc
xrc_wwl_11_21 wwl_11_20 wwl_11_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_21 wbl_10_21 wbl_11_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_21 rwl_11_20 rwl_11_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_21 rbl_10_21 rbl_11_21 rc_unit R0=Rrbl C0=Crbl
xgc_11_22 wwl_11_22 wbl_11_22 rwl_11_22 rbl_11_22 sn_11_22 wos_ros_gc
xrc_wwl_11_22 wwl_11_21 wwl_11_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_22 wbl_10_22 wbl_11_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_22 rwl_11_21 rwl_11_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_22 rbl_10_22 rbl_11_22 rc_unit R0=Rrbl C0=Crbl
xgc_11_23 wwl_11_23 wbl_11_23 rwl_11_23 rbl_11_23 sn_11_23 wos_ros_gc
xrc_wwl_11_23 wwl_11_22 wwl_11_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_23 wbl_10_23 wbl_11_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_23 rwl_11_22 rwl_11_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_23 rbl_10_23 rbl_11_23 rc_unit R0=Rrbl C0=Crbl
xgc_11_24 wwl_11_24 wbl_11_24 rwl_11_24 rbl_11_24 sn_11_24 wos_ros_gc
xrc_wwl_11_24 wwl_11_23 wwl_11_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_24 wbl_10_24 wbl_11_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_24 rwl_11_23 rwl_11_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_24 rbl_10_24 rbl_11_24 rc_unit R0=Rrbl C0=Crbl
xgc_11_25 wwl_11_25 wbl_11_25 rwl_11_25 rbl_11_25 sn_11_25 wos_ros_gc
xrc_wwl_11_25 wwl_11_24 wwl_11_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_25 wbl_10_25 wbl_11_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_25 rwl_11_24 rwl_11_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_25 rbl_10_25 rbl_11_25 rc_unit R0=Rrbl C0=Crbl
xgc_11_26 wwl_11_26 wbl_11_26 rwl_11_26 rbl_11_26 sn_11_26 wos_ros_gc
xrc_wwl_11_26 wwl_11_25 wwl_11_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_26 wbl_10_26 wbl_11_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_26 rwl_11_25 rwl_11_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_26 rbl_10_26 rbl_11_26 rc_unit R0=Rrbl C0=Crbl
xgc_11_27 wwl_11_27 wbl_11_27 rwl_11_27 rbl_11_27 sn_11_27 wos_ros_gc
xrc_wwl_11_27 wwl_11_26 wwl_11_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_27 wbl_10_27 wbl_11_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_27 rwl_11_26 rwl_11_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_27 rbl_10_27 rbl_11_27 rc_unit R0=Rrbl C0=Crbl
xgc_11_28 wwl_11_28 wbl_11_28 rwl_11_28 rbl_11_28 sn_11_28 wos_ros_gc
xrc_wwl_11_28 wwl_11_27 wwl_11_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_28 wbl_10_28 wbl_11_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_28 rwl_11_27 rwl_11_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_28 rbl_10_28 rbl_11_28 rc_unit R0=Rrbl C0=Crbl
xgc_11_29 wwl_11_29 wbl_11_29 rwl_11_29 rbl_11_29 sn_11_29 wos_ros_gc
xrc_wwl_11_29 wwl_11_28 wwl_11_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_29 wbl_10_29 wbl_11_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_29 rwl_11_28 rwl_11_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_29 rbl_10_29 rbl_11_29 rc_unit R0=Rrbl C0=Crbl
xgc_11_30 wwl_11_30 wbl_11_30 rwl_11_30 rbl_11_30 sn_11_30 wos_ros_gc
xrc_wwl_11_30 wwl_11_29 wwl_11_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_30 wbl_10_30 wbl_11_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_30 rwl_11_29 rwl_11_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_30 rbl_10_30 rbl_11_30 rc_unit R0=Rrbl C0=Crbl
xgc_11_31 wwl_11_31 wbl_11_31 rwl_11_31 rbl_11_31 sn_11_31 wos_ros_gc
xrc_wwl_11_31 wwl_11_30 wwl_11_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_11_31 wbl_10_31 wbl_11_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_11_31 rwl_11_30 rwl_11_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_11_31 rbl_10_31 rbl_11_31 rc_unit R0=Rrbl C0=Crbl
xgc_12_0 wwl_12_0 wbl_12_0 rwl_12_0 rbl_12_0 sn_12_0 wos_ros_gc
xrc_wwl_12_0 wwl_12 wwl_12_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_0 wbl_11_0 wbl_12_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_0 rwl_12 rwl_12_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_0 rbl_11_0 rbl_12_0 rc_unit R0=Rrbl C0=Crbl
xgc_12_1 wwl_12_1 wbl_12_1 rwl_12_1 rbl_12_1 sn_12_1 wos_ros_gc
xrc_wwl_12_1 wwl_12_0 wwl_12_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_1 wbl_11_1 wbl_12_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_1 rwl_12_0 rwl_12_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_1 rbl_11_1 rbl_12_1 rc_unit R0=Rrbl C0=Crbl
xgc_12_2 wwl_12_2 wbl_12_2 rwl_12_2 rbl_12_2 sn_12_2 wos_ros_gc
xrc_wwl_12_2 wwl_12_1 wwl_12_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_2 wbl_11_2 wbl_12_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_2 rwl_12_1 rwl_12_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_2 rbl_11_2 rbl_12_2 rc_unit R0=Rrbl C0=Crbl
xgc_12_3 wwl_12_3 wbl_12_3 rwl_12_3 rbl_12_3 sn_12_3 wos_ros_gc
xrc_wwl_12_3 wwl_12_2 wwl_12_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_3 wbl_11_3 wbl_12_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_3 rwl_12_2 rwl_12_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_3 rbl_11_3 rbl_12_3 rc_unit R0=Rrbl C0=Crbl
xgc_12_4 wwl_12_4 wbl_12_4 rwl_12_4 rbl_12_4 sn_12_4 wos_ros_gc
xrc_wwl_12_4 wwl_12_3 wwl_12_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_4 wbl_11_4 wbl_12_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_4 rwl_12_3 rwl_12_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_4 rbl_11_4 rbl_12_4 rc_unit R0=Rrbl C0=Crbl
xgc_12_5 wwl_12_5 wbl_12_5 rwl_12_5 rbl_12_5 sn_12_5 wos_ros_gc
xrc_wwl_12_5 wwl_12_4 wwl_12_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_5 wbl_11_5 wbl_12_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_5 rwl_12_4 rwl_12_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_5 rbl_11_5 rbl_12_5 rc_unit R0=Rrbl C0=Crbl
xgc_12_6 wwl_12_6 wbl_12_6 rwl_12_6 rbl_12_6 sn_12_6 wos_ros_gc
xrc_wwl_12_6 wwl_12_5 wwl_12_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_6 wbl_11_6 wbl_12_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_6 rwl_12_5 rwl_12_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_6 rbl_11_6 rbl_12_6 rc_unit R0=Rrbl C0=Crbl
xgc_12_7 wwl_12_7 wbl_12_7 rwl_12_7 rbl_12_7 sn_12_7 wos_ros_gc
xrc_wwl_12_7 wwl_12_6 wwl_12_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_7 wbl_11_7 wbl_12_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_7 rwl_12_6 rwl_12_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_7 rbl_11_7 rbl_12_7 rc_unit R0=Rrbl C0=Crbl
xgc_12_8 wwl_12_8 wbl_12_8 rwl_12_8 rbl_12_8 sn_12_8 wos_ros_gc
xrc_wwl_12_8 wwl_12_7 wwl_12_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_8 wbl_11_8 wbl_12_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_8 rwl_12_7 rwl_12_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_8 rbl_11_8 rbl_12_8 rc_unit R0=Rrbl C0=Crbl
xgc_12_9 wwl_12_9 wbl_12_9 rwl_12_9 rbl_12_9 sn_12_9 wos_ros_gc
xrc_wwl_12_9 wwl_12_8 wwl_12_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_9 wbl_11_9 wbl_12_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_9 rwl_12_8 rwl_12_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_9 rbl_11_9 rbl_12_9 rc_unit R0=Rrbl C0=Crbl
xgc_12_10 wwl_12_10 wbl_12_10 rwl_12_10 rbl_12_10 sn_12_10 wos_ros_gc
xrc_wwl_12_10 wwl_12_9 wwl_12_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_10 wbl_11_10 wbl_12_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_10 rwl_12_9 rwl_12_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_10 rbl_11_10 rbl_12_10 rc_unit R0=Rrbl C0=Crbl
xgc_12_11 wwl_12_11 wbl_12_11 rwl_12_11 rbl_12_11 sn_12_11 wos_ros_gc
xrc_wwl_12_11 wwl_12_10 wwl_12_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_11 wbl_11_11 wbl_12_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_11 rwl_12_10 rwl_12_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_11 rbl_11_11 rbl_12_11 rc_unit R0=Rrbl C0=Crbl
xgc_12_12 wwl_12_12 wbl_12_12 rwl_12_12 rbl_12_12 sn_12_12 wos_ros_gc
xrc_wwl_12_12 wwl_12_11 wwl_12_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_12 wbl_11_12 wbl_12_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_12 rwl_12_11 rwl_12_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_12 rbl_11_12 rbl_12_12 rc_unit R0=Rrbl C0=Crbl
xgc_12_13 wwl_12_13 wbl_12_13 rwl_12_13 rbl_12_13 sn_12_13 wos_ros_gc
xrc_wwl_12_13 wwl_12_12 wwl_12_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_13 wbl_11_13 wbl_12_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_13 rwl_12_12 rwl_12_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_13 rbl_11_13 rbl_12_13 rc_unit R0=Rrbl C0=Crbl
xgc_12_14 wwl_12_14 wbl_12_14 rwl_12_14 rbl_12_14 sn_12_14 wos_ros_gc
xrc_wwl_12_14 wwl_12_13 wwl_12_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_14 wbl_11_14 wbl_12_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_14 rwl_12_13 rwl_12_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_14 rbl_11_14 rbl_12_14 rc_unit R0=Rrbl C0=Crbl
xgc_12_15 wwl_12_15 wbl_12_15 rwl_12_15 rbl_12_15 sn_12_15 wos_ros_gc
xrc_wwl_12_15 wwl_12_14 wwl_12_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_15 wbl_11_15 wbl_12_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_15 rwl_12_14 rwl_12_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_15 rbl_11_15 rbl_12_15 rc_unit R0=Rrbl C0=Crbl
xgc_12_16 wwl_12_16 wbl_12_16 rwl_12_16 rbl_12_16 sn_12_16 wos_ros_gc
xrc_wwl_12_16 wwl_12_15 wwl_12_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_16 wbl_11_16 wbl_12_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_16 rwl_12_15 rwl_12_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_16 rbl_11_16 rbl_12_16 rc_unit R0=Rrbl C0=Crbl
xgc_12_17 wwl_12_17 wbl_12_17 rwl_12_17 rbl_12_17 sn_12_17 wos_ros_gc
xrc_wwl_12_17 wwl_12_16 wwl_12_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_17 wbl_11_17 wbl_12_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_17 rwl_12_16 rwl_12_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_17 rbl_11_17 rbl_12_17 rc_unit R0=Rrbl C0=Crbl
xgc_12_18 wwl_12_18 wbl_12_18 rwl_12_18 rbl_12_18 sn_12_18 wos_ros_gc
xrc_wwl_12_18 wwl_12_17 wwl_12_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_18 wbl_11_18 wbl_12_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_18 rwl_12_17 rwl_12_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_18 rbl_11_18 rbl_12_18 rc_unit R0=Rrbl C0=Crbl
xgc_12_19 wwl_12_19 wbl_12_19 rwl_12_19 rbl_12_19 sn_12_19 wos_ros_gc
xrc_wwl_12_19 wwl_12_18 wwl_12_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_19 wbl_11_19 wbl_12_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_19 rwl_12_18 rwl_12_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_19 rbl_11_19 rbl_12_19 rc_unit R0=Rrbl C0=Crbl
xgc_12_20 wwl_12_20 wbl_12_20 rwl_12_20 rbl_12_20 sn_12_20 wos_ros_gc
xrc_wwl_12_20 wwl_12_19 wwl_12_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_20 wbl_11_20 wbl_12_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_20 rwl_12_19 rwl_12_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_20 rbl_11_20 rbl_12_20 rc_unit R0=Rrbl C0=Crbl
xgc_12_21 wwl_12_21 wbl_12_21 rwl_12_21 rbl_12_21 sn_12_21 wos_ros_gc
xrc_wwl_12_21 wwl_12_20 wwl_12_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_21 wbl_11_21 wbl_12_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_21 rwl_12_20 rwl_12_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_21 rbl_11_21 rbl_12_21 rc_unit R0=Rrbl C0=Crbl
xgc_12_22 wwl_12_22 wbl_12_22 rwl_12_22 rbl_12_22 sn_12_22 wos_ros_gc
xrc_wwl_12_22 wwl_12_21 wwl_12_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_22 wbl_11_22 wbl_12_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_22 rwl_12_21 rwl_12_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_22 rbl_11_22 rbl_12_22 rc_unit R0=Rrbl C0=Crbl
xgc_12_23 wwl_12_23 wbl_12_23 rwl_12_23 rbl_12_23 sn_12_23 wos_ros_gc
xrc_wwl_12_23 wwl_12_22 wwl_12_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_23 wbl_11_23 wbl_12_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_23 rwl_12_22 rwl_12_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_23 rbl_11_23 rbl_12_23 rc_unit R0=Rrbl C0=Crbl
xgc_12_24 wwl_12_24 wbl_12_24 rwl_12_24 rbl_12_24 sn_12_24 wos_ros_gc
xrc_wwl_12_24 wwl_12_23 wwl_12_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_24 wbl_11_24 wbl_12_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_24 rwl_12_23 rwl_12_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_24 rbl_11_24 rbl_12_24 rc_unit R0=Rrbl C0=Crbl
xgc_12_25 wwl_12_25 wbl_12_25 rwl_12_25 rbl_12_25 sn_12_25 wos_ros_gc
xrc_wwl_12_25 wwl_12_24 wwl_12_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_25 wbl_11_25 wbl_12_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_25 rwl_12_24 rwl_12_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_25 rbl_11_25 rbl_12_25 rc_unit R0=Rrbl C0=Crbl
xgc_12_26 wwl_12_26 wbl_12_26 rwl_12_26 rbl_12_26 sn_12_26 wos_ros_gc
xrc_wwl_12_26 wwl_12_25 wwl_12_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_26 wbl_11_26 wbl_12_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_26 rwl_12_25 rwl_12_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_26 rbl_11_26 rbl_12_26 rc_unit R0=Rrbl C0=Crbl
xgc_12_27 wwl_12_27 wbl_12_27 rwl_12_27 rbl_12_27 sn_12_27 wos_ros_gc
xrc_wwl_12_27 wwl_12_26 wwl_12_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_27 wbl_11_27 wbl_12_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_27 rwl_12_26 rwl_12_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_27 rbl_11_27 rbl_12_27 rc_unit R0=Rrbl C0=Crbl
xgc_12_28 wwl_12_28 wbl_12_28 rwl_12_28 rbl_12_28 sn_12_28 wos_ros_gc
xrc_wwl_12_28 wwl_12_27 wwl_12_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_28 wbl_11_28 wbl_12_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_28 rwl_12_27 rwl_12_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_28 rbl_11_28 rbl_12_28 rc_unit R0=Rrbl C0=Crbl
xgc_12_29 wwl_12_29 wbl_12_29 rwl_12_29 rbl_12_29 sn_12_29 wos_ros_gc
xrc_wwl_12_29 wwl_12_28 wwl_12_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_29 wbl_11_29 wbl_12_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_29 rwl_12_28 rwl_12_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_29 rbl_11_29 rbl_12_29 rc_unit R0=Rrbl C0=Crbl
xgc_12_30 wwl_12_30 wbl_12_30 rwl_12_30 rbl_12_30 sn_12_30 wos_ros_gc
xrc_wwl_12_30 wwl_12_29 wwl_12_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_30 wbl_11_30 wbl_12_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_30 rwl_12_29 rwl_12_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_30 rbl_11_30 rbl_12_30 rc_unit R0=Rrbl C0=Crbl
xgc_12_31 wwl_12_31 wbl_12_31 rwl_12_31 rbl_12_31 sn_12_31 wos_ros_gc
xrc_wwl_12_31 wwl_12_30 wwl_12_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_12_31 wbl_11_31 wbl_12_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_12_31 rwl_12_30 rwl_12_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_12_31 rbl_11_31 rbl_12_31 rc_unit R0=Rrbl C0=Crbl
xgc_13_0 wwl_13_0 wbl_13_0 rwl_13_0 rbl_13_0 sn_13_0 wos_ros_gc
xrc_wwl_13_0 wwl_13 wwl_13_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_0 wbl_12_0 wbl_13_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_0 rwl_13 rwl_13_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_0 rbl_12_0 rbl_13_0 rc_unit R0=Rrbl C0=Crbl
xgc_13_1 wwl_13_1 wbl_13_1 rwl_13_1 rbl_13_1 sn_13_1 wos_ros_gc
xrc_wwl_13_1 wwl_13_0 wwl_13_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_1 wbl_12_1 wbl_13_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_1 rwl_13_0 rwl_13_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_1 rbl_12_1 rbl_13_1 rc_unit R0=Rrbl C0=Crbl
xgc_13_2 wwl_13_2 wbl_13_2 rwl_13_2 rbl_13_2 sn_13_2 wos_ros_gc
xrc_wwl_13_2 wwl_13_1 wwl_13_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_2 wbl_12_2 wbl_13_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_2 rwl_13_1 rwl_13_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_2 rbl_12_2 rbl_13_2 rc_unit R0=Rrbl C0=Crbl
xgc_13_3 wwl_13_3 wbl_13_3 rwl_13_3 rbl_13_3 sn_13_3 wos_ros_gc
xrc_wwl_13_3 wwl_13_2 wwl_13_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_3 wbl_12_3 wbl_13_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_3 rwl_13_2 rwl_13_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_3 rbl_12_3 rbl_13_3 rc_unit R0=Rrbl C0=Crbl
xgc_13_4 wwl_13_4 wbl_13_4 rwl_13_4 rbl_13_4 sn_13_4 wos_ros_gc
xrc_wwl_13_4 wwl_13_3 wwl_13_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_4 wbl_12_4 wbl_13_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_4 rwl_13_3 rwl_13_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_4 rbl_12_4 rbl_13_4 rc_unit R0=Rrbl C0=Crbl
xgc_13_5 wwl_13_5 wbl_13_5 rwl_13_5 rbl_13_5 sn_13_5 wos_ros_gc
xrc_wwl_13_5 wwl_13_4 wwl_13_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_5 wbl_12_5 wbl_13_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_5 rwl_13_4 rwl_13_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_5 rbl_12_5 rbl_13_5 rc_unit R0=Rrbl C0=Crbl
xgc_13_6 wwl_13_6 wbl_13_6 rwl_13_6 rbl_13_6 sn_13_6 wos_ros_gc
xrc_wwl_13_6 wwl_13_5 wwl_13_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_6 wbl_12_6 wbl_13_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_6 rwl_13_5 rwl_13_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_6 rbl_12_6 rbl_13_6 rc_unit R0=Rrbl C0=Crbl
xgc_13_7 wwl_13_7 wbl_13_7 rwl_13_7 rbl_13_7 sn_13_7 wos_ros_gc
xrc_wwl_13_7 wwl_13_6 wwl_13_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_7 wbl_12_7 wbl_13_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_7 rwl_13_6 rwl_13_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_7 rbl_12_7 rbl_13_7 rc_unit R0=Rrbl C0=Crbl
xgc_13_8 wwl_13_8 wbl_13_8 rwl_13_8 rbl_13_8 sn_13_8 wos_ros_gc
xrc_wwl_13_8 wwl_13_7 wwl_13_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_8 wbl_12_8 wbl_13_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_8 rwl_13_7 rwl_13_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_8 rbl_12_8 rbl_13_8 rc_unit R0=Rrbl C0=Crbl
xgc_13_9 wwl_13_9 wbl_13_9 rwl_13_9 rbl_13_9 sn_13_9 wos_ros_gc
xrc_wwl_13_9 wwl_13_8 wwl_13_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_9 wbl_12_9 wbl_13_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_9 rwl_13_8 rwl_13_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_9 rbl_12_9 rbl_13_9 rc_unit R0=Rrbl C0=Crbl
xgc_13_10 wwl_13_10 wbl_13_10 rwl_13_10 rbl_13_10 sn_13_10 wos_ros_gc
xrc_wwl_13_10 wwl_13_9 wwl_13_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_10 wbl_12_10 wbl_13_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_10 rwl_13_9 rwl_13_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_10 rbl_12_10 rbl_13_10 rc_unit R0=Rrbl C0=Crbl
xgc_13_11 wwl_13_11 wbl_13_11 rwl_13_11 rbl_13_11 sn_13_11 wos_ros_gc
xrc_wwl_13_11 wwl_13_10 wwl_13_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_11 wbl_12_11 wbl_13_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_11 rwl_13_10 rwl_13_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_11 rbl_12_11 rbl_13_11 rc_unit R0=Rrbl C0=Crbl
xgc_13_12 wwl_13_12 wbl_13_12 rwl_13_12 rbl_13_12 sn_13_12 wos_ros_gc
xrc_wwl_13_12 wwl_13_11 wwl_13_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_12 wbl_12_12 wbl_13_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_12 rwl_13_11 rwl_13_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_12 rbl_12_12 rbl_13_12 rc_unit R0=Rrbl C0=Crbl
xgc_13_13 wwl_13_13 wbl_13_13 rwl_13_13 rbl_13_13 sn_13_13 wos_ros_gc
xrc_wwl_13_13 wwl_13_12 wwl_13_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_13 wbl_12_13 wbl_13_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_13 rwl_13_12 rwl_13_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_13 rbl_12_13 rbl_13_13 rc_unit R0=Rrbl C0=Crbl
xgc_13_14 wwl_13_14 wbl_13_14 rwl_13_14 rbl_13_14 sn_13_14 wos_ros_gc
xrc_wwl_13_14 wwl_13_13 wwl_13_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_14 wbl_12_14 wbl_13_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_14 rwl_13_13 rwl_13_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_14 rbl_12_14 rbl_13_14 rc_unit R0=Rrbl C0=Crbl
xgc_13_15 wwl_13_15 wbl_13_15 rwl_13_15 rbl_13_15 sn_13_15 wos_ros_gc
xrc_wwl_13_15 wwl_13_14 wwl_13_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_15 wbl_12_15 wbl_13_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_15 rwl_13_14 rwl_13_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_15 rbl_12_15 rbl_13_15 rc_unit R0=Rrbl C0=Crbl
xgc_13_16 wwl_13_16 wbl_13_16 rwl_13_16 rbl_13_16 sn_13_16 wos_ros_gc
xrc_wwl_13_16 wwl_13_15 wwl_13_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_16 wbl_12_16 wbl_13_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_16 rwl_13_15 rwl_13_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_16 rbl_12_16 rbl_13_16 rc_unit R0=Rrbl C0=Crbl
xgc_13_17 wwl_13_17 wbl_13_17 rwl_13_17 rbl_13_17 sn_13_17 wos_ros_gc
xrc_wwl_13_17 wwl_13_16 wwl_13_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_17 wbl_12_17 wbl_13_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_17 rwl_13_16 rwl_13_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_17 rbl_12_17 rbl_13_17 rc_unit R0=Rrbl C0=Crbl
xgc_13_18 wwl_13_18 wbl_13_18 rwl_13_18 rbl_13_18 sn_13_18 wos_ros_gc
xrc_wwl_13_18 wwl_13_17 wwl_13_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_18 wbl_12_18 wbl_13_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_18 rwl_13_17 rwl_13_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_18 rbl_12_18 rbl_13_18 rc_unit R0=Rrbl C0=Crbl
xgc_13_19 wwl_13_19 wbl_13_19 rwl_13_19 rbl_13_19 sn_13_19 wos_ros_gc
xrc_wwl_13_19 wwl_13_18 wwl_13_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_19 wbl_12_19 wbl_13_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_19 rwl_13_18 rwl_13_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_19 rbl_12_19 rbl_13_19 rc_unit R0=Rrbl C0=Crbl
xgc_13_20 wwl_13_20 wbl_13_20 rwl_13_20 rbl_13_20 sn_13_20 wos_ros_gc
xrc_wwl_13_20 wwl_13_19 wwl_13_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_20 wbl_12_20 wbl_13_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_20 rwl_13_19 rwl_13_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_20 rbl_12_20 rbl_13_20 rc_unit R0=Rrbl C0=Crbl
xgc_13_21 wwl_13_21 wbl_13_21 rwl_13_21 rbl_13_21 sn_13_21 wos_ros_gc
xrc_wwl_13_21 wwl_13_20 wwl_13_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_21 wbl_12_21 wbl_13_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_21 rwl_13_20 rwl_13_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_21 rbl_12_21 rbl_13_21 rc_unit R0=Rrbl C0=Crbl
xgc_13_22 wwl_13_22 wbl_13_22 rwl_13_22 rbl_13_22 sn_13_22 wos_ros_gc
xrc_wwl_13_22 wwl_13_21 wwl_13_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_22 wbl_12_22 wbl_13_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_22 rwl_13_21 rwl_13_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_22 rbl_12_22 rbl_13_22 rc_unit R0=Rrbl C0=Crbl
xgc_13_23 wwl_13_23 wbl_13_23 rwl_13_23 rbl_13_23 sn_13_23 wos_ros_gc
xrc_wwl_13_23 wwl_13_22 wwl_13_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_23 wbl_12_23 wbl_13_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_23 rwl_13_22 rwl_13_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_23 rbl_12_23 rbl_13_23 rc_unit R0=Rrbl C0=Crbl
xgc_13_24 wwl_13_24 wbl_13_24 rwl_13_24 rbl_13_24 sn_13_24 wos_ros_gc
xrc_wwl_13_24 wwl_13_23 wwl_13_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_24 wbl_12_24 wbl_13_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_24 rwl_13_23 rwl_13_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_24 rbl_12_24 rbl_13_24 rc_unit R0=Rrbl C0=Crbl
xgc_13_25 wwl_13_25 wbl_13_25 rwl_13_25 rbl_13_25 sn_13_25 wos_ros_gc
xrc_wwl_13_25 wwl_13_24 wwl_13_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_25 wbl_12_25 wbl_13_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_25 rwl_13_24 rwl_13_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_25 rbl_12_25 rbl_13_25 rc_unit R0=Rrbl C0=Crbl
xgc_13_26 wwl_13_26 wbl_13_26 rwl_13_26 rbl_13_26 sn_13_26 wos_ros_gc
xrc_wwl_13_26 wwl_13_25 wwl_13_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_26 wbl_12_26 wbl_13_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_26 rwl_13_25 rwl_13_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_26 rbl_12_26 rbl_13_26 rc_unit R0=Rrbl C0=Crbl
xgc_13_27 wwl_13_27 wbl_13_27 rwl_13_27 rbl_13_27 sn_13_27 wos_ros_gc
xrc_wwl_13_27 wwl_13_26 wwl_13_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_27 wbl_12_27 wbl_13_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_27 rwl_13_26 rwl_13_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_27 rbl_12_27 rbl_13_27 rc_unit R0=Rrbl C0=Crbl
xgc_13_28 wwl_13_28 wbl_13_28 rwl_13_28 rbl_13_28 sn_13_28 wos_ros_gc
xrc_wwl_13_28 wwl_13_27 wwl_13_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_28 wbl_12_28 wbl_13_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_28 rwl_13_27 rwl_13_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_28 rbl_12_28 rbl_13_28 rc_unit R0=Rrbl C0=Crbl
xgc_13_29 wwl_13_29 wbl_13_29 rwl_13_29 rbl_13_29 sn_13_29 wos_ros_gc
xrc_wwl_13_29 wwl_13_28 wwl_13_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_29 wbl_12_29 wbl_13_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_29 rwl_13_28 rwl_13_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_29 rbl_12_29 rbl_13_29 rc_unit R0=Rrbl C0=Crbl
xgc_13_30 wwl_13_30 wbl_13_30 rwl_13_30 rbl_13_30 sn_13_30 wos_ros_gc
xrc_wwl_13_30 wwl_13_29 wwl_13_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_30 wbl_12_30 wbl_13_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_30 rwl_13_29 rwl_13_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_30 rbl_12_30 rbl_13_30 rc_unit R0=Rrbl C0=Crbl
xgc_13_31 wwl_13_31 wbl_13_31 rwl_13_31 rbl_13_31 sn_13_31 wos_ros_gc
xrc_wwl_13_31 wwl_13_30 wwl_13_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_13_31 wbl_12_31 wbl_13_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_13_31 rwl_13_30 rwl_13_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_13_31 rbl_12_31 rbl_13_31 rc_unit R0=Rrbl C0=Crbl
xgc_14_0 wwl_14_0 wbl_14_0 rwl_14_0 rbl_14_0 sn_14_0 wos_ros_gc
xrc_wwl_14_0 wwl_14 wwl_14_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_0 wbl_13_0 wbl_14_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_0 rwl_14 rwl_14_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_0 rbl_13_0 rbl_14_0 rc_unit R0=Rrbl C0=Crbl
xgc_14_1 wwl_14_1 wbl_14_1 rwl_14_1 rbl_14_1 sn_14_1 wos_ros_gc
xrc_wwl_14_1 wwl_14_0 wwl_14_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_1 wbl_13_1 wbl_14_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_1 rwl_14_0 rwl_14_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_1 rbl_13_1 rbl_14_1 rc_unit R0=Rrbl C0=Crbl
xgc_14_2 wwl_14_2 wbl_14_2 rwl_14_2 rbl_14_2 sn_14_2 wos_ros_gc
xrc_wwl_14_2 wwl_14_1 wwl_14_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_2 wbl_13_2 wbl_14_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_2 rwl_14_1 rwl_14_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_2 rbl_13_2 rbl_14_2 rc_unit R0=Rrbl C0=Crbl
xgc_14_3 wwl_14_3 wbl_14_3 rwl_14_3 rbl_14_3 sn_14_3 wos_ros_gc
xrc_wwl_14_3 wwl_14_2 wwl_14_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_3 wbl_13_3 wbl_14_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_3 rwl_14_2 rwl_14_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_3 rbl_13_3 rbl_14_3 rc_unit R0=Rrbl C0=Crbl
xgc_14_4 wwl_14_4 wbl_14_4 rwl_14_4 rbl_14_4 sn_14_4 wos_ros_gc
xrc_wwl_14_4 wwl_14_3 wwl_14_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_4 wbl_13_4 wbl_14_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_4 rwl_14_3 rwl_14_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_4 rbl_13_4 rbl_14_4 rc_unit R0=Rrbl C0=Crbl
xgc_14_5 wwl_14_5 wbl_14_5 rwl_14_5 rbl_14_5 sn_14_5 wos_ros_gc
xrc_wwl_14_5 wwl_14_4 wwl_14_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_5 wbl_13_5 wbl_14_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_5 rwl_14_4 rwl_14_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_5 rbl_13_5 rbl_14_5 rc_unit R0=Rrbl C0=Crbl
xgc_14_6 wwl_14_6 wbl_14_6 rwl_14_6 rbl_14_6 sn_14_6 wos_ros_gc
xrc_wwl_14_6 wwl_14_5 wwl_14_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_6 wbl_13_6 wbl_14_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_6 rwl_14_5 rwl_14_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_6 rbl_13_6 rbl_14_6 rc_unit R0=Rrbl C0=Crbl
xgc_14_7 wwl_14_7 wbl_14_7 rwl_14_7 rbl_14_7 sn_14_7 wos_ros_gc
xrc_wwl_14_7 wwl_14_6 wwl_14_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_7 wbl_13_7 wbl_14_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_7 rwl_14_6 rwl_14_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_7 rbl_13_7 rbl_14_7 rc_unit R0=Rrbl C0=Crbl
xgc_14_8 wwl_14_8 wbl_14_8 rwl_14_8 rbl_14_8 sn_14_8 wos_ros_gc
xrc_wwl_14_8 wwl_14_7 wwl_14_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_8 wbl_13_8 wbl_14_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_8 rwl_14_7 rwl_14_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_8 rbl_13_8 rbl_14_8 rc_unit R0=Rrbl C0=Crbl
xgc_14_9 wwl_14_9 wbl_14_9 rwl_14_9 rbl_14_9 sn_14_9 wos_ros_gc
xrc_wwl_14_9 wwl_14_8 wwl_14_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_9 wbl_13_9 wbl_14_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_9 rwl_14_8 rwl_14_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_9 rbl_13_9 rbl_14_9 rc_unit R0=Rrbl C0=Crbl
xgc_14_10 wwl_14_10 wbl_14_10 rwl_14_10 rbl_14_10 sn_14_10 wos_ros_gc
xrc_wwl_14_10 wwl_14_9 wwl_14_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_10 wbl_13_10 wbl_14_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_10 rwl_14_9 rwl_14_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_10 rbl_13_10 rbl_14_10 rc_unit R0=Rrbl C0=Crbl
xgc_14_11 wwl_14_11 wbl_14_11 rwl_14_11 rbl_14_11 sn_14_11 wos_ros_gc
xrc_wwl_14_11 wwl_14_10 wwl_14_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_11 wbl_13_11 wbl_14_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_11 rwl_14_10 rwl_14_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_11 rbl_13_11 rbl_14_11 rc_unit R0=Rrbl C0=Crbl
xgc_14_12 wwl_14_12 wbl_14_12 rwl_14_12 rbl_14_12 sn_14_12 wos_ros_gc
xrc_wwl_14_12 wwl_14_11 wwl_14_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_12 wbl_13_12 wbl_14_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_12 rwl_14_11 rwl_14_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_12 rbl_13_12 rbl_14_12 rc_unit R0=Rrbl C0=Crbl
xgc_14_13 wwl_14_13 wbl_14_13 rwl_14_13 rbl_14_13 sn_14_13 wos_ros_gc
xrc_wwl_14_13 wwl_14_12 wwl_14_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_13 wbl_13_13 wbl_14_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_13 rwl_14_12 rwl_14_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_13 rbl_13_13 rbl_14_13 rc_unit R0=Rrbl C0=Crbl
xgc_14_14 wwl_14_14 wbl_14_14 rwl_14_14 rbl_14_14 sn_14_14 wos_ros_gc
xrc_wwl_14_14 wwl_14_13 wwl_14_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_14 wbl_13_14 wbl_14_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_14 rwl_14_13 rwl_14_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_14 rbl_13_14 rbl_14_14 rc_unit R0=Rrbl C0=Crbl
xgc_14_15 wwl_14_15 wbl_14_15 rwl_14_15 rbl_14_15 sn_14_15 wos_ros_gc
xrc_wwl_14_15 wwl_14_14 wwl_14_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_15 wbl_13_15 wbl_14_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_15 rwl_14_14 rwl_14_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_15 rbl_13_15 rbl_14_15 rc_unit R0=Rrbl C0=Crbl
xgc_14_16 wwl_14_16 wbl_14_16 rwl_14_16 rbl_14_16 sn_14_16 wos_ros_gc
xrc_wwl_14_16 wwl_14_15 wwl_14_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_16 wbl_13_16 wbl_14_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_16 rwl_14_15 rwl_14_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_16 rbl_13_16 rbl_14_16 rc_unit R0=Rrbl C0=Crbl
xgc_14_17 wwl_14_17 wbl_14_17 rwl_14_17 rbl_14_17 sn_14_17 wos_ros_gc
xrc_wwl_14_17 wwl_14_16 wwl_14_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_17 wbl_13_17 wbl_14_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_17 rwl_14_16 rwl_14_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_17 rbl_13_17 rbl_14_17 rc_unit R0=Rrbl C0=Crbl
xgc_14_18 wwl_14_18 wbl_14_18 rwl_14_18 rbl_14_18 sn_14_18 wos_ros_gc
xrc_wwl_14_18 wwl_14_17 wwl_14_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_18 wbl_13_18 wbl_14_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_18 rwl_14_17 rwl_14_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_18 rbl_13_18 rbl_14_18 rc_unit R0=Rrbl C0=Crbl
xgc_14_19 wwl_14_19 wbl_14_19 rwl_14_19 rbl_14_19 sn_14_19 wos_ros_gc
xrc_wwl_14_19 wwl_14_18 wwl_14_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_19 wbl_13_19 wbl_14_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_19 rwl_14_18 rwl_14_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_19 rbl_13_19 rbl_14_19 rc_unit R0=Rrbl C0=Crbl
xgc_14_20 wwl_14_20 wbl_14_20 rwl_14_20 rbl_14_20 sn_14_20 wos_ros_gc
xrc_wwl_14_20 wwl_14_19 wwl_14_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_20 wbl_13_20 wbl_14_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_20 rwl_14_19 rwl_14_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_20 rbl_13_20 rbl_14_20 rc_unit R0=Rrbl C0=Crbl
xgc_14_21 wwl_14_21 wbl_14_21 rwl_14_21 rbl_14_21 sn_14_21 wos_ros_gc
xrc_wwl_14_21 wwl_14_20 wwl_14_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_21 wbl_13_21 wbl_14_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_21 rwl_14_20 rwl_14_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_21 rbl_13_21 rbl_14_21 rc_unit R0=Rrbl C0=Crbl
xgc_14_22 wwl_14_22 wbl_14_22 rwl_14_22 rbl_14_22 sn_14_22 wos_ros_gc
xrc_wwl_14_22 wwl_14_21 wwl_14_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_22 wbl_13_22 wbl_14_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_22 rwl_14_21 rwl_14_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_22 rbl_13_22 rbl_14_22 rc_unit R0=Rrbl C0=Crbl
xgc_14_23 wwl_14_23 wbl_14_23 rwl_14_23 rbl_14_23 sn_14_23 wos_ros_gc
xrc_wwl_14_23 wwl_14_22 wwl_14_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_23 wbl_13_23 wbl_14_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_23 rwl_14_22 rwl_14_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_23 rbl_13_23 rbl_14_23 rc_unit R0=Rrbl C0=Crbl
xgc_14_24 wwl_14_24 wbl_14_24 rwl_14_24 rbl_14_24 sn_14_24 wos_ros_gc
xrc_wwl_14_24 wwl_14_23 wwl_14_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_24 wbl_13_24 wbl_14_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_24 rwl_14_23 rwl_14_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_24 rbl_13_24 rbl_14_24 rc_unit R0=Rrbl C0=Crbl
xgc_14_25 wwl_14_25 wbl_14_25 rwl_14_25 rbl_14_25 sn_14_25 wos_ros_gc
xrc_wwl_14_25 wwl_14_24 wwl_14_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_25 wbl_13_25 wbl_14_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_25 rwl_14_24 rwl_14_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_25 rbl_13_25 rbl_14_25 rc_unit R0=Rrbl C0=Crbl
xgc_14_26 wwl_14_26 wbl_14_26 rwl_14_26 rbl_14_26 sn_14_26 wos_ros_gc
xrc_wwl_14_26 wwl_14_25 wwl_14_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_26 wbl_13_26 wbl_14_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_26 rwl_14_25 rwl_14_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_26 rbl_13_26 rbl_14_26 rc_unit R0=Rrbl C0=Crbl
xgc_14_27 wwl_14_27 wbl_14_27 rwl_14_27 rbl_14_27 sn_14_27 wos_ros_gc
xrc_wwl_14_27 wwl_14_26 wwl_14_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_27 wbl_13_27 wbl_14_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_27 rwl_14_26 rwl_14_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_27 rbl_13_27 rbl_14_27 rc_unit R0=Rrbl C0=Crbl
xgc_14_28 wwl_14_28 wbl_14_28 rwl_14_28 rbl_14_28 sn_14_28 wos_ros_gc
xrc_wwl_14_28 wwl_14_27 wwl_14_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_28 wbl_13_28 wbl_14_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_28 rwl_14_27 rwl_14_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_28 rbl_13_28 rbl_14_28 rc_unit R0=Rrbl C0=Crbl
xgc_14_29 wwl_14_29 wbl_14_29 rwl_14_29 rbl_14_29 sn_14_29 wos_ros_gc
xrc_wwl_14_29 wwl_14_28 wwl_14_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_29 wbl_13_29 wbl_14_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_29 rwl_14_28 rwl_14_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_29 rbl_13_29 rbl_14_29 rc_unit R0=Rrbl C0=Crbl
xgc_14_30 wwl_14_30 wbl_14_30 rwl_14_30 rbl_14_30 sn_14_30 wos_ros_gc
xrc_wwl_14_30 wwl_14_29 wwl_14_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_30 wbl_13_30 wbl_14_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_30 rwl_14_29 rwl_14_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_30 rbl_13_30 rbl_14_30 rc_unit R0=Rrbl C0=Crbl
xgc_14_31 wwl_14_31 wbl_14_31 rwl_14_31 rbl_14_31 sn_14_31 wos_ros_gc
xrc_wwl_14_31 wwl_14_30 wwl_14_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_14_31 wbl_13_31 wbl_14_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_14_31 rwl_14_30 rwl_14_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_14_31 rbl_13_31 rbl_14_31 rc_unit R0=Rrbl C0=Crbl
xgc_15_0 wwl_15_0 wbl_15_0 rwl_15_0 rbl_15_0 sn_15_0 wos_ros_gc
xrc_wwl_15_0 wwl_15 wwl_15_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_0 wbl_14_0 wbl_15_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_0 rwl_15 rwl_15_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_0 rbl_14_0 rbl_15_0 rc_unit R0=Rrbl C0=Crbl
xgc_15_1 wwl_15_1 wbl_15_1 rwl_15_1 rbl_15_1 sn_15_1 wos_ros_gc
xrc_wwl_15_1 wwl_15_0 wwl_15_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_1 wbl_14_1 wbl_15_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_1 rwl_15_0 rwl_15_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_1 rbl_14_1 rbl_15_1 rc_unit R0=Rrbl C0=Crbl
xgc_15_2 wwl_15_2 wbl_15_2 rwl_15_2 rbl_15_2 sn_15_2 wos_ros_gc
xrc_wwl_15_2 wwl_15_1 wwl_15_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_2 wbl_14_2 wbl_15_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_2 rwl_15_1 rwl_15_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_2 rbl_14_2 rbl_15_2 rc_unit R0=Rrbl C0=Crbl
xgc_15_3 wwl_15_3 wbl_15_3 rwl_15_3 rbl_15_3 sn_15_3 wos_ros_gc
xrc_wwl_15_3 wwl_15_2 wwl_15_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_3 wbl_14_3 wbl_15_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_3 rwl_15_2 rwl_15_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_3 rbl_14_3 rbl_15_3 rc_unit R0=Rrbl C0=Crbl
xgc_15_4 wwl_15_4 wbl_15_4 rwl_15_4 rbl_15_4 sn_15_4 wos_ros_gc
xrc_wwl_15_4 wwl_15_3 wwl_15_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_4 wbl_14_4 wbl_15_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_4 rwl_15_3 rwl_15_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_4 rbl_14_4 rbl_15_4 rc_unit R0=Rrbl C0=Crbl
xgc_15_5 wwl_15_5 wbl_15_5 rwl_15_5 rbl_15_5 sn_15_5 wos_ros_gc
xrc_wwl_15_5 wwl_15_4 wwl_15_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_5 wbl_14_5 wbl_15_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_5 rwl_15_4 rwl_15_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_5 rbl_14_5 rbl_15_5 rc_unit R0=Rrbl C0=Crbl
xgc_15_6 wwl_15_6 wbl_15_6 rwl_15_6 rbl_15_6 sn_15_6 wos_ros_gc
xrc_wwl_15_6 wwl_15_5 wwl_15_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_6 wbl_14_6 wbl_15_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_6 rwl_15_5 rwl_15_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_6 rbl_14_6 rbl_15_6 rc_unit R0=Rrbl C0=Crbl
xgc_15_7 wwl_15_7 wbl_15_7 rwl_15_7 rbl_15_7 sn_15_7 wos_ros_gc
xrc_wwl_15_7 wwl_15_6 wwl_15_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_7 wbl_14_7 wbl_15_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_7 rwl_15_6 rwl_15_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_7 rbl_14_7 rbl_15_7 rc_unit R0=Rrbl C0=Crbl
xgc_15_8 wwl_15_8 wbl_15_8 rwl_15_8 rbl_15_8 sn_15_8 wos_ros_gc
xrc_wwl_15_8 wwl_15_7 wwl_15_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_8 wbl_14_8 wbl_15_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_8 rwl_15_7 rwl_15_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_8 rbl_14_8 rbl_15_8 rc_unit R0=Rrbl C0=Crbl
xgc_15_9 wwl_15_9 wbl_15_9 rwl_15_9 rbl_15_9 sn_15_9 wos_ros_gc
xrc_wwl_15_9 wwl_15_8 wwl_15_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_9 wbl_14_9 wbl_15_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_9 rwl_15_8 rwl_15_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_9 rbl_14_9 rbl_15_9 rc_unit R0=Rrbl C0=Crbl
xgc_15_10 wwl_15_10 wbl_15_10 rwl_15_10 rbl_15_10 sn_15_10 wos_ros_gc
xrc_wwl_15_10 wwl_15_9 wwl_15_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_10 wbl_14_10 wbl_15_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_10 rwl_15_9 rwl_15_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_10 rbl_14_10 rbl_15_10 rc_unit R0=Rrbl C0=Crbl
xgc_15_11 wwl_15_11 wbl_15_11 rwl_15_11 rbl_15_11 sn_15_11 wos_ros_gc
xrc_wwl_15_11 wwl_15_10 wwl_15_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_11 wbl_14_11 wbl_15_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_11 rwl_15_10 rwl_15_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_11 rbl_14_11 rbl_15_11 rc_unit R0=Rrbl C0=Crbl
xgc_15_12 wwl_15_12 wbl_15_12 rwl_15_12 rbl_15_12 sn_15_12 wos_ros_gc
xrc_wwl_15_12 wwl_15_11 wwl_15_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_12 wbl_14_12 wbl_15_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_12 rwl_15_11 rwl_15_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_12 rbl_14_12 rbl_15_12 rc_unit R0=Rrbl C0=Crbl
xgc_15_13 wwl_15_13 wbl_15_13 rwl_15_13 rbl_15_13 sn_15_13 wos_ros_gc
xrc_wwl_15_13 wwl_15_12 wwl_15_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_13 wbl_14_13 wbl_15_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_13 rwl_15_12 rwl_15_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_13 rbl_14_13 rbl_15_13 rc_unit R0=Rrbl C0=Crbl
xgc_15_14 wwl_15_14 wbl_15_14 rwl_15_14 rbl_15_14 sn_15_14 wos_ros_gc
xrc_wwl_15_14 wwl_15_13 wwl_15_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_14 wbl_14_14 wbl_15_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_14 rwl_15_13 rwl_15_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_14 rbl_14_14 rbl_15_14 rc_unit R0=Rrbl C0=Crbl
xgc_15_15 wwl_15_15 wbl_15_15 rwl_15_15 rbl_15_15 sn_15_15 wos_ros_gc
xrc_wwl_15_15 wwl_15_14 wwl_15_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_15 wbl_14_15 wbl_15_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_15 rwl_15_14 rwl_15_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_15 rbl_14_15 rbl_15_15 rc_unit R0=Rrbl C0=Crbl
xgc_15_16 wwl_15_16 wbl_15_16 rwl_15_16 rbl_15_16 sn_15_16 wos_ros_gc
xrc_wwl_15_16 wwl_15_15 wwl_15_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_16 wbl_14_16 wbl_15_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_16 rwl_15_15 rwl_15_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_16 rbl_14_16 rbl_15_16 rc_unit R0=Rrbl C0=Crbl
xgc_15_17 wwl_15_17 wbl_15_17 rwl_15_17 rbl_15_17 sn_15_17 wos_ros_gc
xrc_wwl_15_17 wwl_15_16 wwl_15_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_17 wbl_14_17 wbl_15_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_17 rwl_15_16 rwl_15_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_17 rbl_14_17 rbl_15_17 rc_unit R0=Rrbl C0=Crbl
xgc_15_18 wwl_15_18 wbl_15_18 rwl_15_18 rbl_15_18 sn_15_18 wos_ros_gc
xrc_wwl_15_18 wwl_15_17 wwl_15_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_18 wbl_14_18 wbl_15_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_18 rwl_15_17 rwl_15_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_18 rbl_14_18 rbl_15_18 rc_unit R0=Rrbl C0=Crbl
xgc_15_19 wwl_15_19 wbl_15_19 rwl_15_19 rbl_15_19 sn_15_19 wos_ros_gc
xrc_wwl_15_19 wwl_15_18 wwl_15_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_19 wbl_14_19 wbl_15_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_19 rwl_15_18 rwl_15_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_19 rbl_14_19 rbl_15_19 rc_unit R0=Rrbl C0=Crbl
xgc_15_20 wwl_15_20 wbl_15_20 rwl_15_20 rbl_15_20 sn_15_20 wos_ros_gc
xrc_wwl_15_20 wwl_15_19 wwl_15_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_20 wbl_14_20 wbl_15_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_20 rwl_15_19 rwl_15_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_20 rbl_14_20 rbl_15_20 rc_unit R0=Rrbl C0=Crbl
xgc_15_21 wwl_15_21 wbl_15_21 rwl_15_21 rbl_15_21 sn_15_21 wos_ros_gc
xrc_wwl_15_21 wwl_15_20 wwl_15_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_21 wbl_14_21 wbl_15_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_21 rwl_15_20 rwl_15_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_21 rbl_14_21 rbl_15_21 rc_unit R0=Rrbl C0=Crbl
xgc_15_22 wwl_15_22 wbl_15_22 rwl_15_22 rbl_15_22 sn_15_22 wos_ros_gc
xrc_wwl_15_22 wwl_15_21 wwl_15_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_22 wbl_14_22 wbl_15_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_22 rwl_15_21 rwl_15_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_22 rbl_14_22 rbl_15_22 rc_unit R0=Rrbl C0=Crbl
xgc_15_23 wwl_15_23 wbl_15_23 rwl_15_23 rbl_15_23 sn_15_23 wos_ros_gc
xrc_wwl_15_23 wwl_15_22 wwl_15_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_23 wbl_14_23 wbl_15_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_23 rwl_15_22 rwl_15_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_23 rbl_14_23 rbl_15_23 rc_unit R0=Rrbl C0=Crbl
xgc_15_24 wwl_15_24 wbl_15_24 rwl_15_24 rbl_15_24 sn_15_24 wos_ros_gc
xrc_wwl_15_24 wwl_15_23 wwl_15_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_24 wbl_14_24 wbl_15_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_24 rwl_15_23 rwl_15_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_24 rbl_14_24 rbl_15_24 rc_unit R0=Rrbl C0=Crbl
xgc_15_25 wwl_15_25 wbl_15_25 rwl_15_25 rbl_15_25 sn_15_25 wos_ros_gc
xrc_wwl_15_25 wwl_15_24 wwl_15_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_25 wbl_14_25 wbl_15_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_25 rwl_15_24 rwl_15_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_25 rbl_14_25 rbl_15_25 rc_unit R0=Rrbl C0=Crbl
xgc_15_26 wwl_15_26 wbl_15_26 rwl_15_26 rbl_15_26 sn_15_26 wos_ros_gc
xrc_wwl_15_26 wwl_15_25 wwl_15_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_26 wbl_14_26 wbl_15_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_26 rwl_15_25 rwl_15_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_26 rbl_14_26 rbl_15_26 rc_unit R0=Rrbl C0=Crbl
xgc_15_27 wwl_15_27 wbl_15_27 rwl_15_27 rbl_15_27 sn_15_27 wos_ros_gc
xrc_wwl_15_27 wwl_15_26 wwl_15_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_27 wbl_14_27 wbl_15_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_27 rwl_15_26 rwl_15_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_27 rbl_14_27 rbl_15_27 rc_unit R0=Rrbl C0=Crbl
xgc_15_28 wwl_15_28 wbl_15_28 rwl_15_28 rbl_15_28 sn_15_28 wos_ros_gc
xrc_wwl_15_28 wwl_15_27 wwl_15_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_28 wbl_14_28 wbl_15_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_28 rwl_15_27 rwl_15_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_28 rbl_14_28 rbl_15_28 rc_unit R0=Rrbl C0=Crbl
xgc_15_29 wwl_15_29 wbl_15_29 rwl_15_29 rbl_15_29 sn_15_29 wos_ros_gc
xrc_wwl_15_29 wwl_15_28 wwl_15_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_29 wbl_14_29 wbl_15_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_29 rwl_15_28 rwl_15_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_29 rbl_14_29 rbl_15_29 rc_unit R0=Rrbl C0=Crbl
xgc_15_30 wwl_15_30 wbl_15_30 rwl_15_30 rbl_15_30 sn_15_30 wos_ros_gc
xrc_wwl_15_30 wwl_15_29 wwl_15_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_30 wbl_14_30 wbl_15_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_30 rwl_15_29 rwl_15_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_30 rbl_14_30 rbl_15_30 rc_unit R0=Rrbl C0=Crbl
xgc_15_31 wwl_15_31 wbl_15_31 rwl_15_31 rbl_15_31 sn_15_31 wos_ros_gc
xrc_wwl_15_31 wwl_15_30 wwl_15_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_15_31 wbl_14_31 wbl_15_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_15_31 rwl_15_30 rwl_15_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_15_31 rbl_14_31 rbl_15_31 rc_unit R0=Rrbl C0=Crbl
xgc_16_0 wwl_16_0 wbl_16_0 rwl_16_0 rbl_16_0 sn_16_0 wos_ros_gc
xrc_wwl_16_0 wwl_16 wwl_16_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_0 wbl_15_0 wbl_16_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_0 rwl_16 rwl_16_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_0 rbl_15_0 rbl_16_0 rc_unit R0=Rrbl C0=Crbl
xgc_16_1 wwl_16_1 wbl_16_1 rwl_16_1 rbl_16_1 sn_16_1 wos_ros_gc
xrc_wwl_16_1 wwl_16_0 wwl_16_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_1 wbl_15_1 wbl_16_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_1 rwl_16_0 rwl_16_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_1 rbl_15_1 rbl_16_1 rc_unit R0=Rrbl C0=Crbl
xgc_16_2 wwl_16_2 wbl_16_2 rwl_16_2 rbl_16_2 sn_16_2 wos_ros_gc
xrc_wwl_16_2 wwl_16_1 wwl_16_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_2 wbl_15_2 wbl_16_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_2 rwl_16_1 rwl_16_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_2 rbl_15_2 rbl_16_2 rc_unit R0=Rrbl C0=Crbl
xgc_16_3 wwl_16_3 wbl_16_3 rwl_16_3 rbl_16_3 sn_16_3 wos_ros_gc
xrc_wwl_16_3 wwl_16_2 wwl_16_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_3 wbl_15_3 wbl_16_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_3 rwl_16_2 rwl_16_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_3 rbl_15_3 rbl_16_3 rc_unit R0=Rrbl C0=Crbl
xgc_16_4 wwl_16_4 wbl_16_4 rwl_16_4 rbl_16_4 sn_16_4 wos_ros_gc
xrc_wwl_16_4 wwl_16_3 wwl_16_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_4 wbl_15_4 wbl_16_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_4 rwl_16_3 rwl_16_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_4 rbl_15_4 rbl_16_4 rc_unit R0=Rrbl C0=Crbl
xgc_16_5 wwl_16_5 wbl_16_5 rwl_16_5 rbl_16_5 sn_16_5 wos_ros_gc
xrc_wwl_16_5 wwl_16_4 wwl_16_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_5 wbl_15_5 wbl_16_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_5 rwl_16_4 rwl_16_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_5 rbl_15_5 rbl_16_5 rc_unit R0=Rrbl C0=Crbl
xgc_16_6 wwl_16_6 wbl_16_6 rwl_16_6 rbl_16_6 sn_16_6 wos_ros_gc
xrc_wwl_16_6 wwl_16_5 wwl_16_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_6 wbl_15_6 wbl_16_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_6 rwl_16_5 rwl_16_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_6 rbl_15_6 rbl_16_6 rc_unit R0=Rrbl C0=Crbl
xgc_16_7 wwl_16_7 wbl_16_7 rwl_16_7 rbl_16_7 sn_16_7 wos_ros_gc
xrc_wwl_16_7 wwl_16_6 wwl_16_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_7 wbl_15_7 wbl_16_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_7 rwl_16_6 rwl_16_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_7 rbl_15_7 rbl_16_7 rc_unit R0=Rrbl C0=Crbl
xgc_16_8 wwl_16_8 wbl_16_8 rwl_16_8 rbl_16_8 sn_16_8 wos_ros_gc
xrc_wwl_16_8 wwl_16_7 wwl_16_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_8 wbl_15_8 wbl_16_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_8 rwl_16_7 rwl_16_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_8 rbl_15_8 rbl_16_8 rc_unit R0=Rrbl C0=Crbl
xgc_16_9 wwl_16_9 wbl_16_9 rwl_16_9 rbl_16_9 sn_16_9 wos_ros_gc
xrc_wwl_16_9 wwl_16_8 wwl_16_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_9 wbl_15_9 wbl_16_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_9 rwl_16_8 rwl_16_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_9 rbl_15_9 rbl_16_9 rc_unit R0=Rrbl C0=Crbl
xgc_16_10 wwl_16_10 wbl_16_10 rwl_16_10 rbl_16_10 sn_16_10 wos_ros_gc
xrc_wwl_16_10 wwl_16_9 wwl_16_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_10 wbl_15_10 wbl_16_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_10 rwl_16_9 rwl_16_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_10 rbl_15_10 rbl_16_10 rc_unit R0=Rrbl C0=Crbl
xgc_16_11 wwl_16_11 wbl_16_11 rwl_16_11 rbl_16_11 sn_16_11 wos_ros_gc
xrc_wwl_16_11 wwl_16_10 wwl_16_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_11 wbl_15_11 wbl_16_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_11 rwl_16_10 rwl_16_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_11 rbl_15_11 rbl_16_11 rc_unit R0=Rrbl C0=Crbl
xgc_16_12 wwl_16_12 wbl_16_12 rwl_16_12 rbl_16_12 sn_16_12 wos_ros_gc
xrc_wwl_16_12 wwl_16_11 wwl_16_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_12 wbl_15_12 wbl_16_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_12 rwl_16_11 rwl_16_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_12 rbl_15_12 rbl_16_12 rc_unit R0=Rrbl C0=Crbl
xgc_16_13 wwl_16_13 wbl_16_13 rwl_16_13 rbl_16_13 sn_16_13 wos_ros_gc
xrc_wwl_16_13 wwl_16_12 wwl_16_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_13 wbl_15_13 wbl_16_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_13 rwl_16_12 rwl_16_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_13 rbl_15_13 rbl_16_13 rc_unit R0=Rrbl C0=Crbl
xgc_16_14 wwl_16_14 wbl_16_14 rwl_16_14 rbl_16_14 sn_16_14 wos_ros_gc
xrc_wwl_16_14 wwl_16_13 wwl_16_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_14 wbl_15_14 wbl_16_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_14 rwl_16_13 rwl_16_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_14 rbl_15_14 rbl_16_14 rc_unit R0=Rrbl C0=Crbl
xgc_16_15 wwl_16_15 wbl_16_15 rwl_16_15 rbl_16_15 sn_16_15 wos_ros_gc
xrc_wwl_16_15 wwl_16_14 wwl_16_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_15 wbl_15_15 wbl_16_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_15 rwl_16_14 rwl_16_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_15 rbl_15_15 rbl_16_15 rc_unit R0=Rrbl C0=Crbl
xgc_16_16 wwl_16_16 wbl_16_16 rwl_16_16 rbl_16_16 sn_16_16 wos_ros_gc
xrc_wwl_16_16 wwl_16_15 wwl_16_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_16 wbl_15_16 wbl_16_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_16 rwl_16_15 rwl_16_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_16 rbl_15_16 rbl_16_16 rc_unit R0=Rrbl C0=Crbl
xgc_16_17 wwl_16_17 wbl_16_17 rwl_16_17 rbl_16_17 sn_16_17 wos_ros_gc
xrc_wwl_16_17 wwl_16_16 wwl_16_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_17 wbl_15_17 wbl_16_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_17 rwl_16_16 rwl_16_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_17 rbl_15_17 rbl_16_17 rc_unit R0=Rrbl C0=Crbl
xgc_16_18 wwl_16_18 wbl_16_18 rwl_16_18 rbl_16_18 sn_16_18 wos_ros_gc
xrc_wwl_16_18 wwl_16_17 wwl_16_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_18 wbl_15_18 wbl_16_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_18 rwl_16_17 rwl_16_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_18 rbl_15_18 rbl_16_18 rc_unit R0=Rrbl C0=Crbl
xgc_16_19 wwl_16_19 wbl_16_19 rwl_16_19 rbl_16_19 sn_16_19 wos_ros_gc
xrc_wwl_16_19 wwl_16_18 wwl_16_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_19 wbl_15_19 wbl_16_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_19 rwl_16_18 rwl_16_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_19 rbl_15_19 rbl_16_19 rc_unit R0=Rrbl C0=Crbl
xgc_16_20 wwl_16_20 wbl_16_20 rwl_16_20 rbl_16_20 sn_16_20 wos_ros_gc
xrc_wwl_16_20 wwl_16_19 wwl_16_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_20 wbl_15_20 wbl_16_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_20 rwl_16_19 rwl_16_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_20 rbl_15_20 rbl_16_20 rc_unit R0=Rrbl C0=Crbl
xgc_16_21 wwl_16_21 wbl_16_21 rwl_16_21 rbl_16_21 sn_16_21 wos_ros_gc
xrc_wwl_16_21 wwl_16_20 wwl_16_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_21 wbl_15_21 wbl_16_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_21 rwl_16_20 rwl_16_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_21 rbl_15_21 rbl_16_21 rc_unit R0=Rrbl C0=Crbl
xgc_16_22 wwl_16_22 wbl_16_22 rwl_16_22 rbl_16_22 sn_16_22 wos_ros_gc
xrc_wwl_16_22 wwl_16_21 wwl_16_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_22 wbl_15_22 wbl_16_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_22 rwl_16_21 rwl_16_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_22 rbl_15_22 rbl_16_22 rc_unit R0=Rrbl C0=Crbl
xgc_16_23 wwl_16_23 wbl_16_23 rwl_16_23 rbl_16_23 sn_16_23 wos_ros_gc
xrc_wwl_16_23 wwl_16_22 wwl_16_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_23 wbl_15_23 wbl_16_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_23 rwl_16_22 rwl_16_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_23 rbl_15_23 rbl_16_23 rc_unit R0=Rrbl C0=Crbl
xgc_16_24 wwl_16_24 wbl_16_24 rwl_16_24 rbl_16_24 sn_16_24 wos_ros_gc
xrc_wwl_16_24 wwl_16_23 wwl_16_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_24 wbl_15_24 wbl_16_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_24 rwl_16_23 rwl_16_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_24 rbl_15_24 rbl_16_24 rc_unit R0=Rrbl C0=Crbl
xgc_16_25 wwl_16_25 wbl_16_25 rwl_16_25 rbl_16_25 sn_16_25 wos_ros_gc
xrc_wwl_16_25 wwl_16_24 wwl_16_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_25 wbl_15_25 wbl_16_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_25 rwl_16_24 rwl_16_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_25 rbl_15_25 rbl_16_25 rc_unit R0=Rrbl C0=Crbl
xgc_16_26 wwl_16_26 wbl_16_26 rwl_16_26 rbl_16_26 sn_16_26 wos_ros_gc
xrc_wwl_16_26 wwl_16_25 wwl_16_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_26 wbl_15_26 wbl_16_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_26 rwl_16_25 rwl_16_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_26 rbl_15_26 rbl_16_26 rc_unit R0=Rrbl C0=Crbl
xgc_16_27 wwl_16_27 wbl_16_27 rwl_16_27 rbl_16_27 sn_16_27 wos_ros_gc
xrc_wwl_16_27 wwl_16_26 wwl_16_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_27 wbl_15_27 wbl_16_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_27 rwl_16_26 rwl_16_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_27 rbl_15_27 rbl_16_27 rc_unit R0=Rrbl C0=Crbl
xgc_16_28 wwl_16_28 wbl_16_28 rwl_16_28 rbl_16_28 sn_16_28 wos_ros_gc
xrc_wwl_16_28 wwl_16_27 wwl_16_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_28 wbl_15_28 wbl_16_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_28 rwl_16_27 rwl_16_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_28 rbl_15_28 rbl_16_28 rc_unit R0=Rrbl C0=Crbl
xgc_16_29 wwl_16_29 wbl_16_29 rwl_16_29 rbl_16_29 sn_16_29 wos_ros_gc
xrc_wwl_16_29 wwl_16_28 wwl_16_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_29 wbl_15_29 wbl_16_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_29 rwl_16_28 rwl_16_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_29 rbl_15_29 rbl_16_29 rc_unit R0=Rrbl C0=Crbl
xgc_16_30 wwl_16_30 wbl_16_30 rwl_16_30 rbl_16_30 sn_16_30 wos_ros_gc
xrc_wwl_16_30 wwl_16_29 wwl_16_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_30 wbl_15_30 wbl_16_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_30 rwl_16_29 rwl_16_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_30 rbl_15_30 rbl_16_30 rc_unit R0=Rrbl C0=Crbl
xgc_16_31 wwl_16_31 wbl_16_31 rwl_16_31 rbl_16_31 sn_16_31 wos_ros_gc
xrc_wwl_16_31 wwl_16_30 wwl_16_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_16_31 wbl_15_31 wbl_16_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_16_31 rwl_16_30 rwl_16_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_16_31 rbl_15_31 rbl_16_31 rc_unit R0=Rrbl C0=Crbl
xgc_17_0 wwl_17_0 wbl_17_0 rwl_17_0 rbl_17_0 sn_17_0 wos_ros_gc
xrc_wwl_17_0 wwl_17 wwl_17_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_0 wbl_16_0 wbl_17_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_0 rwl_17 rwl_17_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_0 rbl_16_0 rbl_17_0 rc_unit R0=Rrbl C0=Crbl
xgc_17_1 wwl_17_1 wbl_17_1 rwl_17_1 rbl_17_1 sn_17_1 wos_ros_gc
xrc_wwl_17_1 wwl_17_0 wwl_17_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_1 wbl_16_1 wbl_17_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_1 rwl_17_0 rwl_17_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_1 rbl_16_1 rbl_17_1 rc_unit R0=Rrbl C0=Crbl
xgc_17_2 wwl_17_2 wbl_17_2 rwl_17_2 rbl_17_2 sn_17_2 wos_ros_gc
xrc_wwl_17_2 wwl_17_1 wwl_17_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_2 wbl_16_2 wbl_17_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_2 rwl_17_1 rwl_17_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_2 rbl_16_2 rbl_17_2 rc_unit R0=Rrbl C0=Crbl
xgc_17_3 wwl_17_3 wbl_17_3 rwl_17_3 rbl_17_3 sn_17_3 wos_ros_gc
xrc_wwl_17_3 wwl_17_2 wwl_17_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_3 wbl_16_3 wbl_17_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_3 rwl_17_2 rwl_17_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_3 rbl_16_3 rbl_17_3 rc_unit R0=Rrbl C0=Crbl
xgc_17_4 wwl_17_4 wbl_17_4 rwl_17_4 rbl_17_4 sn_17_4 wos_ros_gc
xrc_wwl_17_4 wwl_17_3 wwl_17_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_4 wbl_16_4 wbl_17_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_4 rwl_17_3 rwl_17_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_4 rbl_16_4 rbl_17_4 rc_unit R0=Rrbl C0=Crbl
xgc_17_5 wwl_17_5 wbl_17_5 rwl_17_5 rbl_17_5 sn_17_5 wos_ros_gc
xrc_wwl_17_5 wwl_17_4 wwl_17_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_5 wbl_16_5 wbl_17_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_5 rwl_17_4 rwl_17_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_5 rbl_16_5 rbl_17_5 rc_unit R0=Rrbl C0=Crbl
xgc_17_6 wwl_17_6 wbl_17_6 rwl_17_6 rbl_17_6 sn_17_6 wos_ros_gc
xrc_wwl_17_6 wwl_17_5 wwl_17_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_6 wbl_16_6 wbl_17_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_6 rwl_17_5 rwl_17_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_6 rbl_16_6 rbl_17_6 rc_unit R0=Rrbl C0=Crbl
xgc_17_7 wwl_17_7 wbl_17_7 rwl_17_7 rbl_17_7 sn_17_7 wos_ros_gc
xrc_wwl_17_7 wwl_17_6 wwl_17_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_7 wbl_16_7 wbl_17_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_7 rwl_17_6 rwl_17_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_7 rbl_16_7 rbl_17_7 rc_unit R0=Rrbl C0=Crbl
xgc_17_8 wwl_17_8 wbl_17_8 rwl_17_8 rbl_17_8 sn_17_8 wos_ros_gc
xrc_wwl_17_8 wwl_17_7 wwl_17_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_8 wbl_16_8 wbl_17_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_8 rwl_17_7 rwl_17_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_8 rbl_16_8 rbl_17_8 rc_unit R0=Rrbl C0=Crbl
xgc_17_9 wwl_17_9 wbl_17_9 rwl_17_9 rbl_17_9 sn_17_9 wos_ros_gc
xrc_wwl_17_9 wwl_17_8 wwl_17_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_9 wbl_16_9 wbl_17_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_9 rwl_17_8 rwl_17_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_9 rbl_16_9 rbl_17_9 rc_unit R0=Rrbl C0=Crbl
xgc_17_10 wwl_17_10 wbl_17_10 rwl_17_10 rbl_17_10 sn_17_10 wos_ros_gc
xrc_wwl_17_10 wwl_17_9 wwl_17_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_10 wbl_16_10 wbl_17_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_10 rwl_17_9 rwl_17_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_10 rbl_16_10 rbl_17_10 rc_unit R0=Rrbl C0=Crbl
xgc_17_11 wwl_17_11 wbl_17_11 rwl_17_11 rbl_17_11 sn_17_11 wos_ros_gc
xrc_wwl_17_11 wwl_17_10 wwl_17_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_11 wbl_16_11 wbl_17_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_11 rwl_17_10 rwl_17_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_11 rbl_16_11 rbl_17_11 rc_unit R0=Rrbl C0=Crbl
xgc_17_12 wwl_17_12 wbl_17_12 rwl_17_12 rbl_17_12 sn_17_12 wos_ros_gc
xrc_wwl_17_12 wwl_17_11 wwl_17_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_12 wbl_16_12 wbl_17_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_12 rwl_17_11 rwl_17_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_12 rbl_16_12 rbl_17_12 rc_unit R0=Rrbl C0=Crbl
xgc_17_13 wwl_17_13 wbl_17_13 rwl_17_13 rbl_17_13 sn_17_13 wos_ros_gc
xrc_wwl_17_13 wwl_17_12 wwl_17_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_13 wbl_16_13 wbl_17_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_13 rwl_17_12 rwl_17_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_13 rbl_16_13 rbl_17_13 rc_unit R0=Rrbl C0=Crbl
xgc_17_14 wwl_17_14 wbl_17_14 rwl_17_14 rbl_17_14 sn_17_14 wos_ros_gc
xrc_wwl_17_14 wwl_17_13 wwl_17_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_14 wbl_16_14 wbl_17_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_14 rwl_17_13 rwl_17_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_14 rbl_16_14 rbl_17_14 rc_unit R0=Rrbl C0=Crbl
xgc_17_15 wwl_17_15 wbl_17_15 rwl_17_15 rbl_17_15 sn_17_15 wos_ros_gc
xrc_wwl_17_15 wwl_17_14 wwl_17_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_15 wbl_16_15 wbl_17_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_15 rwl_17_14 rwl_17_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_15 rbl_16_15 rbl_17_15 rc_unit R0=Rrbl C0=Crbl
xgc_17_16 wwl_17_16 wbl_17_16 rwl_17_16 rbl_17_16 sn_17_16 wos_ros_gc
xrc_wwl_17_16 wwl_17_15 wwl_17_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_16 wbl_16_16 wbl_17_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_16 rwl_17_15 rwl_17_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_16 rbl_16_16 rbl_17_16 rc_unit R0=Rrbl C0=Crbl
xgc_17_17 wwl_17_17 wbl_17_17 rwl_17_17 rbl_17_17 sn_17_17 wos_ros_gc
xrc_wwl_17_17 wwl_17_16 wwl_17_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_17 wbl_16_17 wbl_17_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_17 rwl_17_16 rwl_17_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_17 rbl_16_17 rbl_17_17 rc_unit R0=Rrbl C0=Crbl
xgc_17_18 wwl_17_18 wbl_17_18 rwl_17_18 rbl_17_18 sn_17_18 wos_ros_gc
xrc_wwl_17_18 wwl_17_17 wwl_17_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_18 wbl_16_18 wbl_17_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_18 rwl_17_17 rwl_17_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_18 rbl_16_18 rbl_17_18 rc_unit R0=Rrbl C0=Crbl
xgc_17_19 wwl_17_19 wbl_17_19 rwl_17_19 rbl_17_19 sn_17_19 wos_ros_gc
xrc_wwl_17_19 wwl_17_18 wwl_17_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_19 wbl_16_19 wbl_17_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_19 rwl_17_18 rwl_17_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_19 rbl_16_19 rbl_17_19 rc_unit R0=Rrbl C0=Crbl
xgc_17_20 wwl_17_20 wbl_17_20 rwl_17_20 rbl_17_20 sn_17_20 wos_ros_gc
xrc_wwl_17_20 wwl_17_19 wwl_17_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_20 wbl_16_20 wbl_17_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_20 rwl_17_19 rwl_17_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_20 rbl_16_20 rbl_17_20 rc_unit R0=Rrbl C0=Crbl
xgc_17_21 wwl_17_21 wbl_17_21 rwl_17_21 rbl_17_21 sn_17_21 wos_ros_gc
xrc_wwl_17_21 wwl_17_20 wwl_17_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_21 wbl_16_21 wbl_17_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_21 rwl_17_20 rwl_17_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_21 rbl_16_21 rbl_17_21 rc_unit R0=Rrbl C0=Crbl
xgc_17_22 wwl_17_22 wbl_17_22 rwl_17_22 rbl_17_22 sn_17_22 wos_ros_gc
xrc_wwl_17_22 wwl_17_21 wwl_17_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_22 wbl_16_22 wbl_17_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_22 rwl_17_21 rwl_17_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_22 rbl_16_22 rbl_17_22 rc_unit R0=Rrbl C0=Crbl
xgc_17_23 wwl_17_23 wbl_17_23 rwl_17_23 rbl_17_23 sn_17_23 wos_ros_gc
xrc_wwl_17_23 wwl_17_22 wwl_17_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_23 wbl_16_23 wbl_17_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_23 rwl_17_22 rwl_17_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_23 rbl_16_23 rbl_17_23 rc_unit R0=Rrbl C0=Crbl
xgc_17_24 wwl_17_24 wbl_17_24 rwl_17_24 rbl_17_24 sn_17_24 wos_ros_gc
xrc_wwl_17_24 wwl_17_23 wwl_17_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_24 wbl_16_24 wbl_17_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_24 rwl_17_23 rwl_17_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_24 rbl_16_24 rbl_17_24 rc_unit R0=Rrbl C0=Crbl
xgc_17_25 wwl_17_25 wbl_17_25 rwl_17_25 rbl_17_25 sn_17_25 wos_ros_gc
xrc_wwl_17_25 wwl_17_24 wwl_17_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_25 wbl_16_25 wbl_17_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_25 rwl_17_24 rwl_17_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_25 rbl_16_25 rbl_17_25 rc_unit R0=Rrbl C0=Crbl
xgc_17_26 wwl_17_26 wbl_17_26 rwl_17_26 rbl_17_26 sn_17_26 wos_ros_gc
xrc_wwl_17_26 wwl_17_25 wwl_17_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_26 wbl_16_26 wbl_17_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_26 rwl_17_25 rwl_17_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_26 rbl_16_26 rbl_17_26 rc_unit R0=Rrbl C0=Crbl
xgc_17_27 wwl_17_27 wbl_17_27 rwl_17_27 rbl_17_27 sn_17_27 wos_ros_gc
xrc_wwl_17_27 wwl_17_26 wwl_17_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_27 wbl_16_27 wbl_17_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_27 rwl_17_26 rwl_17_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_27 rbl_16_27 rbl_17_27 rc_unit R0=Rrbl C0=Crbl
xgc_17_28 wwl_17_28 wbl_17_28 rwl_17_28 rbl_17_28 sn_17_28 wos_ros_gc
xrc_wwl_17_28 wwl_17_27 wwl_17_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_28 wbl_16_28 wbl_17_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_28 rwl_17_27 rwl_17_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_28 rbl_16_28 rbl_17_28 rc_unit R0=Rrbl C0=Crbl
xgc_17_29 wwl_17_29 wbl_17_29 rwl_17_29 rbl_17_29 sn_17_29 wos_ros_gc
xrc_wwl_17_29 wwl_17_28 wwl_17_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_29 wbl_16_29 wbl_17_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_29 rwl_17_28 rwl_17_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_29 rbl_16_29 rbl_17_29 rc_unit R0=Rrbl C0=Crbl
xgc_17_30 wwl_17_30 wbl_17_30 rwl_17_30 rbl_17_30 sn_17_30 wos_ros_gc
xrc_wwl_17_30 wwl_17_29 wwl_17_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_30 wbl_16_30 wbl_17_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_30 rwl_17_29 rwl_17_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_30 rbl_16_30 rbl_17_30 rc_unit R0=Rrbl C0=Crbl
xgc_17_31 wwl_17_31 wbl_17_31 rwl_17_31 rbl_17_31 sn_17_31 wos_ros_gc
xrc_wwl_17_31 wwl_17_30 wwl_17_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_17_31 wbl_16_31 wbl_17_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_17_31 rwl_17_30 rwl_17_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_17_31 rbl_16_31 rbl_17_31 rc_unit R0=Rrbl C0=Crbl
xgc_18_0 wwl_18_0 wbl_18_0 rwl_18_0 rbl_18_0 sn_18_0 wos_ros_gc
xrc_wwl_18_0 wwl_18 wwl_18_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_0 wbl_17_0 wbl_18_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_0 rwl_18 rwl_18_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_0 rbl_17_0 rbl_18_0 rc_unit R0=Rrbl C0=Crbl
xgc_18_1 wwl_18_1 wbl_18_1 rwl_18_1 rbl_18_1 sn_18_1 wos_ros_gc
xrc_wwl_18_1 wwl_18_0 wwl_18_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_1 wbl_17_1 wbl_18_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_1 rwl_18_0 rwl_18_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_1 rbl_17_1 rbl_18_1 rc_unit R0=Rrbl C0=Crbl
xgc_18_2 wwl_18_2 wbl_18_2 rwl_18_2 rbl_18_2 sn_18_2 wos_ros_gc
xrc_wwl_18_2 wwl_18_1 wwl_18_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_2 wbl_17_2 wbl_18_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_2 rwl_18_1 rwl_18_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_2 rbl_17_2 rbl_18_2 rc_unit R0=Rrbl C0=Crbl
xgc_18_3 wwl_18_3 wbl_18_3 rwl_18_3 rbl_18_3 sn_18_3 wos_ros_gc
xrc_wwl_18_3 wwl_18_2 wwl_18_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_3 wbl_17_3 wbl_18_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_3 rwl_18_2 rwl_18_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_3 rbl_17_3 rbl_18_3 rc_unit R0=Rrbl C0=Crbl
xgc_18_4 wwl_18_4 wbl_18_4 rwl_18_4 rbl_18_4 sn_18_4 wos_ros_gc
xrc_wwl_18_4 wwl_18_3 wwl_18_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_4 wbl_17_4 wbl_18_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_4 rwl_18_3 rwl_18_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_4 rbl_17_4 rbl_18_4 rc_unit R0=Rrbl C0=Crbl
xgc_18_5 wwl_18_5 wbl_18_5 rwl_18_5 rbl_18_5 sn_18_5 wos_ros_gc
xrc_wwl_18_5 wwl_18_4 wwl_18_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_5 wbl_17_5 wbl_18_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_5 rwl_18_4 rwl_18_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_5 rbl_17_5 rbl_18_5 rc_unit R0=Rrbl C0=Crbl
xgc_18_6 wwl_18_6 wbl_18_6 rwl_18_6 rbl_18_6 sn_18_6 wos_ros_gc
xrc_wwl_18_6 wwl_18_5 wwl_18_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_6 wbl_17_6 wbl_18_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_6 rwl_18_5 rwl_18_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_6 rbl_17_6 rbl_18_6 rc_unit R0=Rrbl C0=Crbl
xgc_18_7 wwl_18_7 wbl_18_7 rwl_18_7 rbl_18_7 sn_18_7 wos_ros_gc
xrc_wwl_18_7 wwl_18_6 wwl_18_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_7 wbl_17_7 wbl_18_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_7 rwl_18_6 rwl_18_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_7 rbl_17_7 rbl_18_7 rc_unit R0=Rrbl C0=Crbl
xgc_18_8 wwl_18_8 wbl_18_8 rwl_18_8 rbl_18_8 sn_18_8 wos_ros_gc
xrc_wwl_18_8 wwl_18_7 wwl_18_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_8 wbl_17_8 wbl_18_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_8 rwl_18_7 rwl_18_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_8 rbl_17_8 rbl_18_8 rc_unit R0=Rrbl C0=Crbl
xgc_18_9 wwl_18_9 wbl_18_9 rwl_18_9 rbl_18_9 sn_18_9 wos_ros_gc
xrc_wwl_18_9 wwl_18_8 wwl_18_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_9 wbl_17_9 wbl_18_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_9 rwl_18_8 rwl_18_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_9 rbl_17_9 rbl_18_9 rc_unit R0=Rrbl C0=Crbl
xgc_18_10 wwl_18_10 wbl_18_10 rwl_18_10 rbl_18_10 sn_18_10 wos_ros_gc
xrc_wwl_18_10 wwl_18_9 wwl_18_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_10 wbl_17_10 wbl_18_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_10 rwl_18_9 rwl_18_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_10 rbl_17_10 rbl_18_10 rc_unit R0=Rrbl C0=Crbl
xgc_18_11 wwl_18_11 wbl_18_11 rwl_18_11 rbl_18_11 sn_18_11 wos_ros_gc
xrc_wwl_18_11 wwl_18_10 wwl_18_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_11 wbl_17_11 wbl_18_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_11 rwl_18_10 rwl_18_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_11 rbl_17_11 rbl_18_11 rc_unit R0=Rrbl C0=Crbl
xgc_18_12 wwl_18_12 wbl_18_12 rwl_18_12 rbl_18_12 sn_18_12 wos_ros_gc
xrc_wwl_18_12 wwl_18_11 wwl_18_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_12 wbl_17_12 wbl_18_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_12 rwl_18_11 rwl_18_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_12 rbl_17_12 rbl_18_12 rc_unit R0=Rrbl C0=Crbl
xgc_18_13 wwl_18_13 wbl_18_13 rwl_18_13 rbl_18_13 sn_18_13 wos_ros_gc
xrc_wwl_18_13 wwl_18_12 wwl_18_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_13 wbl_17_13 wbl_18_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_13 rwl_18_12 rwl_18_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_13 rbl_17_13 rbl_18_13 rc_unit R0=Rrbl C0=Crbl
xgc_18_14 wwl_18_14 wbl_18_14 rwl_18_14 rbl_18_14 sn_18_14 wos_ros_gc
xrc_wwl_18_14 wwl_18_13 wwl_18_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_14 wbl_17_14 wbl_18_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_14 rwl_18_13 rwl_18_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_14 rbl_17_14 rbl_18_14 rc_unit R0=Rrbl C0=Crbl
xgc_18_15 wwl_18_15 wbl_18_15 rwl_18_15 rbl_18_15 sn_18_15 wos_ros_gc
xrc_wwl_18_15 wwl_18_14 wwl_18_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_15 wbl_17_15 wbl_18_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_15 rwl_18_14 rwl_18_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_15 rbl_17_15 rbl_18_15 rc_unit R0=Rrbl C0=Crbl
xgc_18_16 wwl_18_16 wbl_18_16 rwl_18_16 rbl_18_16 sn_18_16 wos_ros_gc
xrc_wwl_18_16 wwl_18_15 wwl_18_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_16 wbl_17_16 wbl_18_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_16 rwl_18_15 rwl_18_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_16 rbl_17_16 rbl_18_16 rc_unit R0=Rrbl C0=Crbl
xgc_18_17 wwl_18_17 wbl_18_17 rwl_18_17 rbl_18_17 sn_18_17 wos_ros_gc
xrc_wwl_18_17 wwl_18_16 wwl_18_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_17 wbl_17_17 wbl_18_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_17 rwl_18_16 rwl_18_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_17 rbl_17_17 rbl_18_17 rc_unit R0=Rrbl C0=Crbl
xgc_18_18 wwl_18_18 wbl_18_18 rwl_18_18 rbl_18_18 sn_18_18 wos_ros_gc
xrc_wwl_18_18 wwl_18_17 wwl_18_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_18 wbl_17_18 wbl_18_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_18 rwl_18_17 rwl_18_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_18 rbl_17_18 rbl_18_18 rc_unit R0=Rrbl C0=Crbl
xgc_18_19 wwl_18_19 wbl_18_19 rwl_18_19 rbl_18_19 sn_18_19 wos_ros_gc
xrc_wwl_18_19 wwl_18_18 wwl_18_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_19 wbl_17_19 wbl_18_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_19 rwl_18_18 rwl_18_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_19 rbl_17_19 rbl_18_19 rc_unit R0=Rrbl C0=Crbl
xgc_18_20 wwl_18_20 wbl_18_20 rwl_18_20 rbl_18_20 sn_18_20 wos_ros_gc
xrc_wwl_18_20 wwl_18_19 wwl_18_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_20 wbl_17_20 wbl_18_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_20 rwl_18_19 rwl_18_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_20 rbl_17_20 rbl_18_20 rc_unit R0=Rrbl C0=Crbl
xgc_18_21 wwl_18_21 wbl_18_21 rwl_18_21 rbl_18_21 sn_18_21 wos_ros_gc
xrc_wwl_18_21 wwl_18_20 wwl_18_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_21 wbl_17_21 wbl_18_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_21 rwl_18_20 rwl_18_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_21 rbl_17_21 rbl_18_21 rc_unit R0=Rrbl C0=Crbl
xgc_18_22 wwl_18_22 wbl_18_22 rwl_18_22 rbl_18_22 sn_18_22 wos_ros_gc
xrc_wwl_18_22 wwl_18_21 wwl_18_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_22 wbl_17_22 wbl_18_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_22 rwl_18_21 rwl_18_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_22 rbl_17_22 rbl_18_22 rc_unit R0=Rrbl C0=Crbl
xgc_18_23 wwl_18_23 wbl_18_23 rwl_18_23 rbl_18_23 sn_18_23 wos_ros_gc
xrc_wwl_18_23 wwl_18_22 wwl_18_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_23 wbl_17_23 wbl_18_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_23 rwl_18_22 rwl_18_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_23 rbl_17_23 rbl_18_23 rc_unit R0=Rrbl C0=Crbl
xgc_18_24 wwl_18_24 wbl_18_24 rwl_18_24 rbl_18_24 sn_18_24 wos_ros_gc
xrc_wwl_18_24 wwl_18_23 wwl_18_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_24 wbl_17_24 wbl_18_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_24 rwl_18_23 rwl_18_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_24 rbl_17_24 rbl_18_24 rc_unit R0=Rrbl C0=Crbl
xgc_18_25 wwl_18_25 wbl_18_25 rwl_18_25 rbl_18_25 sn_18_25 wos_ros_gc
xrc_wwl_18_25 wwl_18_24 wwl_18_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_25 wbl_17_25 wbl_18_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_25 rwl_18_24 rwl_18_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_25 rbl_17_25 rbl_18_25 rc_unit R0=Rrbl C0=Crbl
xgc_18_26 wwl_18_26 wbl_18_26 rwl_18_26 rbl_18_26 sn_18_26 wos_ros_gc
xrc_wwl_18_26 wwl_18_25 wwl_18_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_26 wbl_17_26 wbl_18_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_26 rwl_18_25 rwl_18_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_26 rbl_17_26 rbl_18_26 rc_unit R0=Rrbl C0=Crbl
xgc_18_27 wwl_18_27 wbl_18_27 rwl_18_27 rbl_18_27 sn_18_27 wos_ros_gc
xrc_wwl_18_27 wwl_18_26 wwl_18_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_27 wbl_17_27 wbl_18_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_27 rwl_18_26 rwl_18_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_27 rbl_17_27 rbl_18_27 rc_unit R0=Rrbl C0=Crbl
xgc_18_28 wwl_18_28 wbl_18_28 rwl_18_28 rbl_18_28 sn_18_28 wos_ros_gc
xrc_wwl_18_28 wwl_18_27 wwl_18_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_28 wbl_17_28 wbl_18_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_28 rwl_18_27 rwl_18_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_28 rbl_17_28 rbl_18_28 rc_unit R0=Rrbl C0=Crbl
xgc_18_29 wwl_18_29 wbl_18_29 rwl_18_29 rbl_18_29 sn_18_29 wos_ros_gc
xrc_wwl_18_29 wwl_18_28 wwl_18_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_29 wbl_17_29 wbl_18_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_29 rwl_18_28 rwl_18_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_29 rbl_17_29 rbl_18_29 rc_unit R0=Rrbl C0=Crbl
xgc_18_30 wwl_18_30 wbl_18_30 rwl_18_30 rbl_18_30 sn_18_30 wos_ros_gc
xrc_wwl_18_30 wwl_18_29 wwl_18_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_30 wbl_17_30 wbl_18_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_30 rwl_18_29 rwl_18_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_30 rbl_17_30 rbl_18_30 rc_unit R0=Rrbl C0=Crbl
xgc_18_31 wwl_18_31 wbl_18_31 rwl_18_31 rbl_18_31 sn_18_31 wos_ros_gc
xrc_wwl_18_31 wwl_18_30 wwl_18_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_18_31 wbl_17_31 wbl_18_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_18_31 rwl_18_30 rwl_18_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_18_31 rbl_17_31 rbl_18_31 rc_unit R0=Rrbl C0=Crbl
xgc_19_0 wwl_19_0 wbl_19_0 rwl_19_0 rbl_19_0 sn_19_0 wos_ros_gc
xrc_wwl_19_0 wwl_19 wwl_19_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_0 wbl_18_0 wbl_19_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_0 rwl_19 rwl_19_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_0 rbl_18_0 rbl_19_0 rc_unit R0=Rrbl C0=Crbl
xgc_19_1 wwl_19_1 wbl_19_1 rwl_19_1 rbl_19_1 sn_19_1 wos_ros_gc
xrc_wwl_19_1 wwl_19_0 wwl_19_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_1 wbl_18_1 wbl_19_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_1 rwl_19_0 rwl_19_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_1 rbl_18_1 rbl_19_1 rc_unit R0=Rrbl C0=Crbl
xgc_19_2 wwl_19_2 wbl_19_2 rwl_19_2 rbl_19_2 sn_19_2 wos_ros_gc
xrc_wwl_19_2 wwl_19_1 wwl_19_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_2 wbl_18_2 wbl_19_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_2 rwl_19_1 rwl_19_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_2 rbl_18_2 rbl_19_2 rc_unit R0=Rrbl C0=Crbl
xgc_19_3 wwl_19_3 wbl_19_3 rwl_19_3 rbl_19_3 sn_19_3 wos_ros_gc
xrc_wwl_19_3 wwl_19_2 wwl_19_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_3 wbl_18_3 wbl_19_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_3 rwl_19_2 rwl_19_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_3 rbl_18_3 rbl_19_3 rc_unit R0=Rrbl C0=Crbl
xgc_19_4 wwl_19_4 wbl_19_4 rwl_19_4 rbl_19_4 sn_19_4 wos_ros_gc
xrc_wwl_19_4 wwl_19_3 wwl_19_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_4 wbl_18_4 wbl_19_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_4 rwl_19_3 rwl_19_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_4 rbl_18_4 rbl_19_4 rc_unit R0=Rrbl C0=Crbl
xgc_19_5 wwl_19_5 wbl_19_5 rwl_19_5 rbl_19_5 sn_19_5 wos_ros_gc
xrc_wwl_19_5 wwl_19_4 wwl_19_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_5 wbl_18_5 wbl_19_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_5 rwl_19_4 rwl_19_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_5 rbl_18_5 rbl_19_5 rc_unit R0=Rrbl C0=Crbl
xgc_19_6 wwl_19_6 wbl_19_6 rwl_19_6 rbl_19_6 sn_19_6 wos_ros_gc
xrc_wwl_19_6 wwl_19_5 wwl_19_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_6 wbl_18_6 wbl_19_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_6 rwl_19_5 rwl_19_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_6 rbl_18_6 rbl_19_6 rc_unit R0=Rrbl C0=Crbl
xgc_19_7 wwl_19_7 wbl_19_7 rwl_19_7 rbl_19_7 sn_19_7 wos_ros_gc
xrc_wwl_19_7 wwl_19_6 wwl_19_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_7 wbl_18_7 wbl_19_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_7 rwl_19_6 rwl_19_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_7 rbl_18_7 rbl_19_7 rc_unit R0=Rrbl C0=Crbl
xgc_19_8 wwl_19_8 wbl_19_8 rwl_19_8 rbl_19_8 sn_19_8 wos_ros_gc
xrc_wwl_19_8 wwl_19_7 wwl_19_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_8 wbl_18_8 wbl_19_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_8 rwl_19_7 rwl_19_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_8 rbl_18_8 rbl_19_8 rc_unit R0=Rrbl C0=Crbl
xgc_19_9 wwl_19_9 wbl_19_9 rwl_19_9 rbl_19_9 sn_19_9 wos_ros_gc
xrc_wwl_19_9 wwl_19_8 wwl_19_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_9 wbl_18_9 wbl_19_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_9 rwl_19_8 rwl_19_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_9 rbl_18_9 rbl_19_9 rc_unit R0=Rrbl C0=Crbl
xgc_19_10 wwl_19_10 wbl_19_10 rwl_19_10 rbl_19_10 sn_19_10 wos_ros_gc
xrc_wwl_19_10 wwl_19_9 wwl_19_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_10 wbl_18_10 wbl_19_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_10 rwl_19_9 rwl_19_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_10 rbl_18_10 rbl_19_10 rc_unit R0=Rrbl C0=Crbl
xgc_19_11 wwl_19_11 wbl_19_11 rwl_19_11 rbl_19_11 sn_19_11 wos_ros_gc
xrc_wwl_19_11 wwl_19_10 wwl_19_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_11 wbl_18_11 wbl_19_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_11 rwl_19_10 rwl_19_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_11 rbl_18_11 rbl_19_11 rc_unit R0=Rrbl C0=Crbl
xgc_19_12 wwl_19_12 wbl_19_12 rwl_19_12 rbl_19_12 sn_19_12 wos_ros_gc
xrc_wwl_19_12 wwl_19_11 wwl_19_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_12 wbl_18_12 wbl_19_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_12 rwl_19_11 rwl_19_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_12 rbl_18_12 rbl_19_12 rc_unit R0=Rrbl C0=Crbl
xgc_19_13 wwl_19_13 wbl_19_13 rwl_19_13 rbl_19_13 sn_19_13 wos_ros_gc
xrc_wwl_19_13 wwl_19_12 wwl_19_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_13 wbl_18_13 wbl_19_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_13 rwl_19_12 rwl_19_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_13 rbl_18_13 rbl_19_13 rc_unit R0=Rrbl C0=Crbl
xgc_19_14 wwl_19_14 wbl_19_14 rwl_19_14 rbl_19_14 sn_19_14 wos_ros_gc
xrc_wwl_19_14 wwl_19_13 wwl_19_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_14 wbl_18_14 wbl_19_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_14 rwl_19_13 rwl_19_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_14 rbl_18_14 rbl_19_14 rc_unit R0=Rrbl C0=Crbl
xgc_19_15 wwl_19_15 wbl_19_15 rwl_19_15 rbl_19_15 sn_19_15 wos_ros_gc
xrc_wwl_19_15 wwl_19_14 wwl_19_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_15 wbl_18_15 wbl_19_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_15 rwl_19_14 rwl_19_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_15 rbl_18_15 rbl_19_15 rc_unit R0=Rrbl C0=Crbl
xgc_19_16 wwl_19_16 wbl_19_16 rwl_19_16 rbl_19_16 sn_19_16 wos_ros_gc
xrc_wwl_19_16 wwl_19_15 wwl_19_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_16 wbl_18_16 wbl_19_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_16 rwl_19_15 rwl_19_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_16 rbl_18_16 rbl_19_16 rc_unit R0=Rrbl C0=Crbl
xgc_19_17 wwl_19_17 wbl_19_17 rwl_19_17 rbl_19_17 sn_19_17 wos_ros_gc
xrc_wwl_19_17 wwl_19_16 wwl_19_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_17 wbl_18_17 wbl_19_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_17 rwl_19_16 rwl_19_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_17 rbl_18_17 rbl_19_17 rc_unit R0=Rrbl C0=Crbl
xgc_19_18 wwl_19_18 wbl_19_18 rwl_19_18 rbl_19_18 sn_19_18 wos_ros_gc
xrc_wwl_19_18 wwl_19_17 wwl_19_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_18 wbl_18_18 wbl_19_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_18 rwl_19_17 rwl_19_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_18 rbl_18_18 rbl_19_18 rc_unit R0=Rrbl C0=Crbl
xgc_19_19 wwl_19_19 wbl_19_19 rwl_19_19 rbl_19_19 sn_19_19 wos_ros_gc
xrc_wwl_19_19 wwl_19_18 wwl_19_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_19 wbl_18_19 wbl_19_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_19 rwl_19_18 rwl_19_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_19 rbl_18_19 rbl_19_19 rc_unit R0=Rrbl C0=Crbl
xgc_19_20 wwl_19_20 wbl_19_20 rwl_19_20 rbl_19_20 sn_19_20 wos_ros_gc
xrc_wwl_19_20 wwl_19_19 wwl_19_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_20 wbl_18_20 wbl_19_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_20 rwl_19_19 rwl_19_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_20 rbl_18_20 rbl_19_20 rc_unit R0=Rrbl C0=Crbl
xgc_19_21 wwl_19_21 wbl_19_21 rwl_19_21 rbl_19_21 sn_19_21 wos_ros_gc
xrc_wwl_19_21 wwl_19_20 wwl_19_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_21 wbl_18_21 wbl_19_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_21 rwl_19_20 rwl_19_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_21 rbl_18_21 rbl_19_21 rc_unit R0=Rrbl C0=Crbl
xgc_19_22 wwl_19_22 wbl_19_22 rwl_19_22 rbl_19_22 sn_19_22 wos_ros_gc
xrc_wwl_19_22 wwl_19_21 wwl_19_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_22 wbl_18_22 wbl_19_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_22 rwl_19_21 rwl_19_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_22 rbl_18_22 rbl_19_22 rc_unit R0=Rrbl C0=Crbl
xgc_19_23 wwl_19_23 wbl_19_23 rwl_19_23 rbl_19_23 sn_19_23 wos_ros_gc
xrc_wwl_19_23 wwl_19_22 wwl_19_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_23 wbl_18_23 wbl_19_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_23 rwl_19_22 rwl_19_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_23 rbl_18_23 rbl_19_23 rc_unit R0=Rrbl C0=Crbl
xgc_19_24 wwl_19_24 wbl_19_24 rwl_19_24 rbl_19_24 sn_19_24 wos_ros_gc
xrc_wwl_19_24 wwl_19_23 wwl_19_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_24 wbl_18_24 wbl_19_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_24 rwl_19_23 rwl_19_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_24 rbl_18_24 rbl_19_24 rc_unit R0=Rrbl C0=Crbl
xgc_19_25 wwl_19_25 wbl_19_25 rwl_19_25 rbl_19_25 sn_19_25 wos_ros_gc
xrc_wwl_19_25 wwl_19_24 wwl_19_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_25 wbl_18_25 wbl_19_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_25 rwl_19_24 rwl_19_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_25 rbl_18_25 rbl_19_25 rc_unit R0=Rrbl C0=Crbl
xgc_19_26 wwl_19_26 wbl_19_26 rwl_19_26 rbl_19_26 sn_19_26 wos_ros_gc
xrc_wwl_19_26 wwl_19_25 wwl_19_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_26 wbl_18_26 wbl_19_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_26 rwl_19_25 rwl_19_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_26 rbl_18_26 rbl_19_26 rc_unit R0=Rrbl C0=Crbl
xgc_19_27 wwl_19_27 wbl_19_27 rwl_19_27 rbl_19_27 sn_19_27 wos_ros_gc
xrc_wwl_19_27 wwl_19_26 wwl_19_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_27 wbl_18_27 wbl_19_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_27 rwl_19_26 rwl_19_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_27 rbl_18_27 rbl_19_27 rc_unit R0=Rrbl C0=Crbl
xgc_19_28 wwl_19_28 wbl_19_28 rwl_19_28 rbl_19_28 sn_19_28 wos_ros_gc
xrc_wwl_19_28 wwl_19_27 wwl_19_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_28 wbl_18_28 wbl_19_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_28 rwl_19_27 rwl_19_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_28 rbl_18_28 rbl_19_28 rc_unit R0=Rrbl C0=Crbl
xgc_19_29 wwl_19_29 wbl_19_29 rwl_19_29 rbl_19_29 sn_19_29 wos_ros_gc
xrc_wwl_19_29 wwl_19_28 wwl_19_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_29 wbl_18_29 wbl_19_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_29 rwl_19_28 rwl_19_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_29 rbl_18_29 rbl_19_29 rc_unit R0=Rrbl C0=Crbl
xgc_19_30 wwl_19_30 wbl_19_30 rwl_19_30 rbl_19_30 sn_19_30 wos_ros_gc
xrc_wwl_19_30 wwl_19_29 wwl_19_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_30 wbl_18_30 wbl_19_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_30 rwl_19_29 rwl_19_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_30 rbl_18_30 rbl_19_30 rc_unit R0=Rrbl C0=Crbl
xgc_19_31 wwl_19_31 wbl_19_31 rwl_19_31 rbl_19_31 sn_19_31 wos_ros_gc
xrc_wwl_19_31 wwl_19_30 wwl_19_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_19_31 wbl_18_31 wbl_19_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_19_31 rwl_19_30 rwl_19_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_19_31 rbl_18_31 rbl_19_31 rc_unit R0=Rrbl C0=Crbl
xgc_20_0 wwl_20_0 wbl_20_0 rwl_20_0 rbl_20_0 sn_20_0 wos_ros_gc
xrc_wwl_20_0 wwl_20 wwl_20_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_0 wbl_19_0 wbl_20_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_0 rwl_20 rwl_20_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_0 rbl_19_0 rbl_20_0 rc_unit R0=Rrbl C0=Crbl
xgc_20_1 wwl_20_1 wbl_20_1 rwl_20_1 rbl_20_1 sn_20_1 wos_ros_gc
xrc_wwl_20_1 wwl_20_0 wwl_20_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_1 wbl_19_1 wbl_20_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_1 rwl_20_0 rwl_20_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_1 rbl_19_1 rbl_20_1 rc_unit R0=Rrbl C0=Crbl
xgc_20_2 wwl_20_2 wbl_20_2 rwl_20_2 rbl_20_2 sn_20_2 wos_ros_gc
xrc_wwl_20_2 wwl_20_1 wwl_20_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_2 wbl_19_2 wbl_20_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_2 rwl_20_1 rwl_20_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_2 rbl_19_2 rbl_20_2 rc_unit R0=Rrbl C0=Crbl
xgc_20_3 wwl_20_3 wbl_20_3 rwl_20_3 rbl_20_3 sn_20_3 wos_ros_gc
xrc_wwl_20_3 wwl_20_2 wwl_20_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_3 wbl_19_3 wbl_20_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_3 rwl_20_2 rwl_20_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_3 rbl_19_3 rbl_20_3 rc_unit R0=Rrbl C0=Crbl
xgc_20_4 wwl_20_4 wbl_20_4 rwl_20_4 rbl_20_4 sn_20_4 wos_ros_gc
xrc_wwl_20_4 wwl_20_3 wwl_20_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_4 wbl_19_4 wbl_20_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_4 rwl_20_3 rwl_20_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_4 rbl_19_4 rbl_20_4 rc_unit R0=Rrbl C0=Crbl
xgc_20_5 wwl_20_5 wbl_20_5 rwl_20_5 rbl_20_5 sn_20_5 wos_ros_gc
xrc_wwl_20_5 wwl_20_4 wwl_20_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_5 wbl_19_5 wbl_20_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_5 rwl_20_4 rwl_20_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_5 rbl_19_5 rbl_20_5 rc_unit R0=Rrbl C0=Crbl
xgc_20_6 wwl_20_6 wbl_20_6 rwl_20_6 rbl_20_6 sn_20_6 wos_ros_gc
xrc_wwl_20_6 wwl_20_5 wwl_20_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_6 wbl_19_6 wbl_20_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_6 rwl_20_5 rwl_20_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_6 rbl_19_6 rbl_20_6 rc_unit R0=Rrbl C0=Crbl
xgc_20_7 wwl_20_7 wbl_20_7 rwl_20_7 rbl_20_7 sn_20_7 wos_ros_gc
xrc_wwl_20_7 wwl_20_6 wwl_20_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_7 wbl_19_7 wbl_20_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_7 rwl_20_6 rwl_20_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_7 rbl_19_7 rbl_20_7 rc_unit R0=Rrbl C0=Crbl
xgc_20_8 wwl_20_8 wbl_20_8 rwl_20_8 rbl_20_8 sn_20_8 wos_ros_gc
xrc_wwl_20_8 wwl_20_7 wwl_20_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_8 wbl_19_8 wbl_20_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_8 rwl_20_7 rwl_20_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_8 rbl_19_8 rbl_20_8 rc_unit R0=Rrbl C0=Crbl
xgc_20_9 wwl_20_9 wbl_20_9 rwl_20_9 rbl_20_9 sn_20_9 wos_ros_gc
xrc_wwl_20_9 wwl_20_8 wwl_20_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_9 wbl_19_9 wbl_20_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_9 rwl_20_8 rwl_20_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_9 rbl_19_9 rbl_20_9 rc_unit R0=Rrbl C0=Crbl
xgc_20_10 wwl_20_10 wbl_20_10 rwl_20_10 rbl_20_10 sn_20_10 wos_ros_gc
xrc_wwl_20_10 wwl_20_9 wwl_20_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_10 wbl_19_10 wbl_20_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_10 rwl_20_9 rwl_20_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_10 rbl_19_10 rbl_20_10 rc_unit R0=Rrbl C0=Crbl
xgc_20_11 wwl_20_11 wbl_20_11 rwl_20_11 rbl_20_11 sn_20_11 wos_ros_gc
xrc_wwl_20_11 wwl_20_10 wwl_20_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_11 wbl_19_11 wbl_20_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_11 rwl_20_10 rwl_20_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_11 rbl_19_11 rbl_20_11 rc_unit R0=Rrbl C0=Crbl
xgc_20_12 wwl_20_12 wbl_20_12 rwl_20_12 rbl_20_12 sn_20_12 wos_ros_gc
xrc_wwl_20_12 wwl_20_11 wwl_20_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_12 wbl_19_12 wbl_20_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_12 rwl_20_11 rwl_20_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_12 rbl_19_12 rbl_20_12 rc_unit R0=Rrbl C0=Crbl
xgc_20_13 wwl_20_13 wbl_20_13 rwl_20_13 rbl_20_13 sn_20_13 wos_ros_gc
xrc_wwl_20_13 wwl_20_12 wwl_20_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_13 wbl_19_13 wbl_20_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_13 rwl_20_12 rwl_20_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_13 rbl_19_13 rbl_20_13 rc_unit R0=Rrbl C0=Crbl
xgc_20_14 wwl_20_14 wbl_20_14 rwl_20_14 rbl_20_14 sn_20_14 wos_ros_gc
xrc_wwl_20_14 wwl_20_13 wwl_20_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_14 wbl_19_14 wbl_20_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_14 rwl_20_13 rwl_20_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_14 rbl_19_14 rbl_20_14 rc_unit R0=Rrbl C0=Crbl
xgc_20_15 wwl_20_15 wbl_20_15 rwl_20_15 rbl_20_15 sn_20_15 wos_ros_gc
xrc_wwl_20_15 wwl_20_14 wwl_20_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_15 wbl_19_15 wbl_20_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_15 rwl_20_14 rwl_20_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_15 rbl_19_15 rbl_20_15 rc_unit R0=Rrbl C0=Crbl
xgc_20_16 wwl_20_16 wbl_20_16 rwl_20_16 rbl_20_16 sn_20_16 wos_ros_gc
xrc_wwl_20_16 wwl_20_15 wwl_20_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_16 wbl_19_16 wbl_20_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_16 rwl_20_15 rwl_20_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_16 rbl_19_16 rbl_20_16 rc_unit R0=Rrbl C0=Crbl
xgc_20_17 wwl_20_17 wbl_20_17 rwl_20_17 rbl_20_17 sn_20_17 wos_ros_gc
xrc_wwl_20_17 wwl_20_16 wwl_20_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_17 wbl_19_17 wbl_20_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_17 rwl_20_16 rwl_20_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_17 rbl_19_17 rbl_20_17 rc_unit R0=Rrbl C0=Crbl
xgc_20_18 wwl_20_18 wbl_20_18 rwl_20_18 rbl_20_18 sn_20_18 wos_ros_gc
xrc_wwl_20_18 wwl_20_17 wwl_20_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_18 wbl_19_18 wbl_20_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_18 rwl_20_17 rwl_20_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_18 rbl_19_18 rbl_20_18 rc_unit R0=Rrbl C0=Crbl
xgc_20_19 wwl_20_19 wbl_20_19 rwl_20_19 rbl_20_19 sn_20_19 wos_ros_gc
xrc_wwl_20_19 wwl_20_18 wwl_20_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_19 wbl_19_19 wbl_20_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_19 rwl_20_18 rwl_20_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_19 rbl_19_19 rbl_20_19 rc_unit R0=Rrbl C0=Crbl
xgc_20_20 wwl_20_20 wbl_20_20 rwl_20_20 rbl_20_20 sn_20_20 wos_ros_gc
xrc_wwl_20_20 wwl_20_19 wwl_20_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_20 wbl_19_20 wbl_20_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_20 rwl_20_19 rwl_20_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_20 rbl_19_20 rbl_20_20 rc_unit R0=Rrbl C0=Crbl
xgc_20_21 wwl_20_21 wbl_20_21 rwl_20_21 rbl_20_21 sn_20_21 wos_ros_gc
xrc_wwl_20_21 wwl_20_20 wwl_20_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_21 wbl_19_21 wbl_20_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_21 rwl_20_20 rwl_20_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_21 rbl_19_21 rbl_20_21 rc_unit R0=Rrbl C0=Crbl
xgc_20_22 wwl_20_22 wbl_20_22 rwl_20_22 rbl_20_22 sn_20_22 wos_ros_gc
xrc_wwl_20_22 wwl_20_21 wwl_20_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_22 wbl_19_22 wbl_20_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_22 rwl_20_21 rwl_20_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_22 rbl_19_22 rbl_20_22 rc_unit R0=Rrbl C0=Crbl
xgc_20_23 wwl_20_23 wbl_20_23 rwl_20_23 rbl_20_23 sn_20_23 wos_ros_gc
xrc_wwl_20_23 wwl_20_22 wwl_20_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_23 wbl_19_23 wbl_20_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_23 rwl_20_22 rwl_20_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_23 rbl_19_23 rbl_20_23 rc_unit R0=Rrbl C0=Crbl
xgc_20_24 wwl_20_24 wbl_20_24 rwl_20_24 rbl_20_24 sn_20_24 wos_ros_gc
xrc_wwl_20_24 wwl_20_23 wwl_20_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_24 wbl_19_24 wbl_20_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_24 rwl_20_23 rwl_20_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_24 rbl_19_24 rbl_20_24 rc_unit R0=Rrbl C0=Crbl
xgc_20_25 wwl_20_25 wbl_20_25 rwl_20_25 rbl_20_25 sn_20_25 wos_ros_gc
xrc_wwl_20_25 wwl_20_24 wwl_20_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_25 wbl_19_25 wbl_20_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_25 rwl_20_24 rwl_20_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_25 rbl_19_25 rbl_20_25 rc_unit R0=Rrbl C0=Crbl
xgc_20_26 wwl_20_26 wbl_20_26 rwl_20_26 rbl_20_26 sn_20_26 wos_ros_gc
xrc_wwl_20_26 wwl_20_25 wwl_20_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_26 wbl_19_26 wbl_20_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_26 rwl_20_25 rwl_20_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_26 rbl_19_26 rbl_20_26 rc_unit R0=Rrbl C0=Crbl
xgc_20_27 wwl_20_27 wbl_20_27 rwl_20_27 rbl_20_27 sn_20_27 wos_ros_gc
xrc_wwl_20_27 wwl_20_26 wwl_20_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_27 wbl_19_27 wbl_20_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_27 rwl_20_26 rwl_20_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_27 rbl_19_27 rbl_20_27 rc_unit R0=Rrbl C0=Crbl
xgc_20_28 wwl_20_28 wbl_20_28 rwl_20_28 rbl_20_28 sn_20_28 wos_ros_gc
xrc_wwl_20_28 wwl_20_27 wwl_20_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_28 wbl_19_28 wbl_20_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_28 rwl_20_27 rwl_20_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_28 rbl_19_28 rbl_20_28 rc_unit R0=Rrbl C0=Crbl
xgc_20_29 wwl_20_29 wbl_20_29 rwl_20_29 rbl_20_29 sn_20_29 wos_ros_gc
xrc_wwl_20_29 wwl_20_28 wwl_20_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_29 wbl_19_29 wbl_20_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_29 rwl_20_28 rwl_20_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_29 rbl_19_29 rbl_20_29 rc_unit R0=Rrbl C0=Crbl
xgc_20_30 wwl_20_30 wbl_20_30 rwl_20_30 rbl_20_30 sn_20_30 wos_ros_gc
xrc_wwl_20_30 wwl_20_29 wwl_20_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_30 wbl_19_30 wbl_20_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_30 rwl_20_29 rwl_20_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_30 rbl_19_30 rbl_20_30 rc_unit R0=Rrbl C0=Crbl
xgc_20_31 wwl_20_31 wbl_20_31 rwl_20_31 rbl_20_31 sn_20_31 wos_ros_gc
xrc_wwl_20_31 wwl_20_30 wwl_20_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_20_31 wbl_19_31 wbl_20_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_20_31 rwl_20_30 rwl_20_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_20_31 rbl_19_31 rbl_20_31 rc_unit R0=Rrbl C0=Crbl
xgc_21_0 wwl_21_0 wbl_21_0 rwl_21_0 rbl_21_0 sn_21_0 wos_ros_gc
xrc_wwl_21_0 wwl_21 wwl_21_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_0 wbl_20_0 wbl_21_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_0 rwl_21 rwl_21_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_0 rbl_20_0 rbl_21_0 rc_unit R0=Rrbl C0=Crbl
xgc_21_1 wwl_21_1 wbl_21_1 rwl_21_1 rbl_21_1 sn_21_1 wos_ros_gc
xrc_wwl_21_1 wwl_21_0 wwl_21_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_1 wbl_20_1 wbl_21_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_1 rwl_21_0 rwl_21_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_1 rbl_20_1 rbl_21_1 rc_unit R0=Rrbl C0=Crbl
xgc_21_2 wwl_21_2 wbl_21_2 rwl_21_2 rbl_21_2 sn_21_2 wos_ros_gc
xrc_wwl_21_2 wwl_21_1 wwl_21_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_2 wbl_20_2 wbl_21_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_2 rwl_21_1 rwl_21_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_2 rbl_20_2 rbl_21_2 rc_unit R0=Rrbl C0=Crbl
xgc_21_3 wwl_21_3 wbl_21_3 rwl_21_3 rbl_21_3 sn_21_3 wos_ros_gc
xrc_wwl_21_3 wwl_21_2 wwl_21_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_3 wbl_20_3 wbl_21_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_3 rwl_21_2 rwl_21_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_3 rbl_20_3 rbl_21_3 rc_unit R0=Rrbl C0=Crbl
xgc_21_4 wwl_21_4 wbl_21_4 rwl_21_4 rbl_21_4 sn_21_4 wos_ros_gc
xrc_wwl_21_4 wwl_21_3 wwl_21_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_4 wbl_20_4 wbl_21_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_4 rwl_21_3 rwl_21_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_4 rbl_20_4 rbl_21_4 rc_unit R0=Rrbl C0=Crbl
xgc_21_5 wwl_21_5 wbl_21_5 rwl_21_5 rbl_21_5 sn_21_5 wos_ros_gc
xrc_wwl_21_5 wwl_21_4 wwl_21_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_5 wbl_20_5 wbl_21_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_5 rwl_21_4 rwl_21_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_5 rbl_20_5 rbl_21_5 rc_unit R0=Rrbl C0=Crbl
xgc_21_6 wwl_21_6 wbl_21_6 rwl_21_6 rbl_21_6 sn_21_6 wos_ros_gc
xrc_wwl_21_6 wwl_21_5 wwl_21_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_6 wbl_20_6 wbl_21_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_6 rwl_21_5 rwl_21_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_6 rbl_20_6 rbl_21_6 rc_unit R0=Rrbl C0=Crbl
xgc_21_7 wwl_21_7 wbl_21_7 rwl_21_7 rbl_21_7 sn_21_7 wos_ros_gc
xrc_wwl_21_7 wwl_21_6 wwl_21_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_7 wbl_20_7 wbl_21_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_7 rwl_21_6 rwl_21_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_7 rbl_20_7 rbl_21_7 rc_unit R0=Rrbl C0=Crbl
xgc_21_8 wwl_21_8 wbl_21_8 rwl_21_8 rbl_21_8 sn_21_8 wos_ros_gc
xrc_wwl_21_8 wwl_21_7 wwl_21_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_8 wbl_20_8 wbl_21_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_8 rwl_21_7 rwl_21_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_8 rbl_20_8 rbl_21_8 rc_unit R0=Rrbl C0=Crbl
xgc_21_9 wwl_21_9 wbl_21_9 rwl_21_9 rbl_21_9 sn_21_9 wos_ros_gc
xrc_wwl_21_9 wwl_21_8 wwl_21_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_9 wbl_20_9 wbl_21_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_9 rwl_21_8 rwl_21_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_9 rbl_20_9 rbl_21_9 rc_unit R0=Rrbl C0=Crbl
xgc_21_10 wwl_21_10 wbl_21_10 rwl_21_10 rbl_21_10 sn_21_10 wos_ros_gc
xrc_wwl_21_10 wwl_21_9 wwl_21_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_10 wbl_20_10 wbl_21_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_10 rwl_21_9 rwl_21_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_10 rbl_20_10 rbl_21_10 rc_unit R0=Rrbl C0=Crbl
xgc_21_11 wwl_21_11 wbl_21_11 rwl_21_11 rbl_21_11 sn_21_11 wos_ros_gc
xrc_wwl_21_11 wwl_21_10 wwl_21_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_11 wbl_20_11 wbl_21_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_11 rwl_21_10 rwl_21_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_11 rbl_20_11 rbl_21_11 rc_unit R0=Rrbl C0=Crbl
xgc_21_12 wwl_21_12 wbl_21_12 rwl_21_12 rbl_21_12 sn_21_12 wos_ros_gc
xrc_wwl_21_12 wwl_21_11 wwl_21_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_12 wbl_20_12 wbl_21_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_12 rwl_21_11 rwl_21_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_12 rbl_20_12 rbl_21_12 rc_unit R0=Rrbl C0=Crbl
xgc_21_13 wwl_21_13 wbl_21_13 rwl_21_13 rbl_21_13 sn_21_13 wos_ros_gc
xrc_wwl_21_13 wwl_21_12 wwl_21_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_13 wbl_20_13 wbl_21_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_13 rwl_21_12 rwl_21_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_13 rbl_20_13 rbl_21_13 rc_unit R0=Rrbl C0=Crbl
xgc_21_14 wwl_21_14 wbl_21_14 rwl_21_14 rbl_21_14 sn_21_14 wos_ros_gc
xrc_wwl_21_14 wwl_21_13 wwl_21_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_14 wbl_20_14 wbl_21_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_14 rwl_21_13 rwl_21_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_14 rbl_20_14 rbl_21_14 rc_unit R0=Rrbl C0=Crbl
xgc_21_15 wwl_21_15 wbl_21_15 rwl_21_15 rbl_21_15 sn_21_15 wos_ros_gc
xrc_wwl_21_15 wwl_21_14 wwl_21_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_15 wbl_20_15 wbl_21_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_15 rwl_21_14 rwl_21_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_15 rbl_20_15 rbl_21_15 rc_unit R0=Rrbl C0=Crbl
xgc_21_16 wwl_21_16 wbl_21_16 rwl_21_16 rbl_21_16 sn_21_16 wos_ros_gc
xrc_wwl_21_16 wwl_21_15 wwl_21_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_16 wbl_20_16 wbl_21_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_16 rwl_21_15 rwl_21_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_16 rbl_20_16 rbl_21_16 rc_unit R0=Rrbl C0=Crbl
xgc_21_17 wwl_21_17 wbl_21_17 rwl_21_17 rbl_21_17 sn_21_17 wos_ros_gc
xrc_wwl_21_17 wwl_21_16 wwl_21_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_17 wbl_20_17 wbl_21_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_17 rwl_21_16 rwl_21_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_17 rbl_20_17 rbl_21_17 rc_unit R0=Rrbl C0=Crbl
xgc_21_18 wwl_21_18 wbl_21_18 rwl_21_18 rbl_21_18 sn_21_18 wos_ros_gc
xrc_wwl_21_18 wwl_21_17 wwl_21_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_18 wbl_20_18 wbl_21_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_18 rwl_21_17 rwl_21_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_18 rbl_20_18 rbl_21_18 rc_unit R0=Rrbl C0=Crbl
xgc_21_19 wwl_21_19 wbl_21_19 rwl_21_19 rbl_21_19 sn_21_19 wos_ros_gc
xrc_wwl_21_19 wwl_21_18 wwl_21_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_19 wbl_20_19 wbl_21_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_19 rwl_21_18 rwl_21_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_19 rbl_20_19 rbl_21_19 rc_unit R0=Rrbl C0=Crbl
xgc_21_20 wwl_21_20 wbl_21_20 rwl_21_20 rbl_21_20 sn_21_20 wos_ros_gc
xrc_wwl_21_20 wwl_21_19 wwl_21_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_20 wbl_20_20 wbl_21_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_20 rwl_21_19 rwl_21_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_20 rbl_20_20 rbl_21_20 rc_unit R0=Rrbl C0=Crbl
xgc_21_21 wwl_21_21 wbl_21_21 rwl_21_21 rbl_21_21 sn_21_21 wos_ros_gc
xrc_wwl_21_21 wwl_21_20 wwl_21_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_21 wbl_20_21 wbl_21_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_21 rwl_21_20 rwl_21_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_21 rbl_20_21 rbl_21_21 rc_unit R0=Rrbl C0=Crbl
xgc_21_22 wwl_21_22 wbl_21_22 rwl_21_22 rbl_21_22 sn_21_22 wos_ros_gc
xrc_wwl_21_22 wwl_21_21 wwl_21_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_22 wbl_20_22 wbl_21_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_22 rwl_21_21 rwl_21_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_22 rbl_20_22 rbl_21_22 rc_unit R0=Rrbl C0=Crbl
xgc_21_23 wwl_21_23 wbl_21_23 rwl_21_23 rbl_21_23 sn_21_23 wos_ros_gc
xrc_wwl_21_23 wwl_21_22 wwl_21_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_23 wbl_20_23 wbl_21_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_23 rwl_21_22 rwl_21_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_23 rbl_20_23 rbl_21_23 rc_unit R0=Rrbl C0=Crbl
xgc_21_24 wwl_21_24 wbl_21_24 rwl_21_24 rbl_21_24 sn_21_24 wos_ros_gc
xrc_wwl_21_24 wwl_21_23 wwl_21_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_24 wbl_20_24 wbl_21_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_24 rwl_21_23 rwl_21_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_24 rbl_20_24 rbl_21_24 rc_unit R0=Rrbl C0=Crbl
xgc_21_25 wwl_21_25 wbl_21_25 rwl_21_25 rbl_21_25 sn_21_25 wos_ros_gc
xrc_wwl_21_25 wwl_21_24 wwl_21_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_25 wbl_20_25 wbl_21_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_25 rwl_21_24 rwl_21_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_25 rbl_20_25 rbl_21_25 rc_unit R0=Rrbl C0=Crbl
xgc_21_26 wwl_21_26 wbl_21_26 rwl_21_26 rbl_21_26 sn_21_26 wos_ros_gc
xrc_wwl_21_26 wwl_21_25 wwl_21_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_26 wbl_20_26 wbl_21_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_26 rwl_21_25 rwl_21_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_26 rbl_20_26 rbl_21_26 rc_unit R0=Rrbl C0=Crbl
xgc_21_27 wwl_21_27 wbl_21_27 rwl_21_27 rbl_21_27 sn_21_27 wos_ros_gc
xrc_wwl_21_27 wwl_21_26 wwl_21_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_27 wbl_20_27 wbl_21_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_27 rwl_21_26 rwl_21_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_27 rbl_20_27 rbl_21_27 rc_unit R0=Rrbl C0=Crbl
xgc_21_28 wwl_21_28 wbl_21_28 rwl_21_28 rbl_21_28 sn_21_28 wos_ros_gc
xrc_wwl_21_28 wwl_21_27 wwl_21_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_28 wbl_20_28 wbl_21_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_28 rwl_21_27 rwl_21_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_28 rbl_20_28 rbl_21_28 rc_unit R0=Rrbl C0=Crbl
xgc_21_29 wwl_21_29 wbl_21_29 rwl_21_29 rbl_21_29 sn_21_29 wos_ros_gc
xrc_wwl_21_29 wwl_21_28 wwl_21_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_29 wbl_20_29 wbl_21_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_29 rwl_21_28 rwl_21_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_29 rbl_20_29 rbl_21_29 rc_unit R0=Rrbl C0=Crbl
xgc_21_30 wwl_21_30 wbl_21_30 rwl_21_30 rbl_21_30 sn_21_30 wos_ros_gc
xrc_wwl_21_30 wwl_21_29 wwl_21_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_30 wbl_20_30 wbl_21_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_30 rwl_21_29 rwl_21_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_30 rbl_20_30 rbl_21_30 rc_unit R0=Rrbl C0=Crbl
xgc_21_31 wwl_21_31 wbl_21_31 rwl_21_31 rbl_21_31 sn_21_31 wos_ros_gc
xrc_wwl_21_31 wwl_21_30 wwl_21_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_21_31 wbl_20_31 wbl_21_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_21_31 rwl_21_30 rwl_21_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_21_31 rbl_20_31 rbl_21_31 rc_unit R0=Rrbl C0=Crbl
xgc_22_0 wwl_22_0 wbl_22_0 rwl_22_0 rbl_22_0 sn_22_0 wos_ros_gc
xrc_wwl_22_0 wwl_22 wwl_22_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_0 wbl_21_0 wbl_22_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_0 rwl_22 rwl_22_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_0 rbl_21_0 rbl_22_0 rc_unit R0=Rrbl C0=Crbl
xgc_22_1 wwl_22_1 wbl_22_1 rwl_22_1 rbl_22_1 sn_22_1 wos_ros_gc
xrc_wwl_22_1 wwl_22_0 wwl_22_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_1 wbl_21_1 wbl_22_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_1 rwl_22_0 rwl_22_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_1 rbl_21_1 rbl_22_1 rc_unit R0=Rrbl C0=Crbl
xgc_22_2 wwl_22_2 wbl_22_2 rwl_22_2 rbl_22_2 sn_22_2 wos_ros_gc
xrc_wwl_22_2 wwl_22_1 wwl_22_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_2 wbl_21_2 wbl_22_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_2 rwl_22_1 rwl_22_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_2 rbl_21_2 rbl_22_2 rc_unit R0=Rrbl C0=Crbl
xgc_22_3 wwl_22_3 wbl_22_3 rwl_22_3 rbl_22_3 sn_22_3 wos_ros_gc
xrc_wwl_22_3 wwl_22_2 wwl_22_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_3 wbl_21_3 wbl_22_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_3 rwl_22_2 rwl_22_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_3 rbl_21_3 rbl_22_3 rc_unit R0=Rrbl C0=Crbl
xgc_22_4 wwl_22_4 wbl_22_4 rwl_22_4 rbl_22_4 sn_22_4 wos_ros_gc
xrc_wwl_22_4 wwl_22_3 wwl_22_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_4 wbl_21_4 wbl_22_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_4 rwl_22_3 rwl_22_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_4 rbl_21_4 rbl_22_4 rc_unit R0=Rrbl C0=Crbl
xgc_22_5 wwl_22_5 wbl_22_5 rwl_22_5 rbl_22_5 sn_22_5 wos_ros_gc
xrc_wwl_22_5 wwl_22_4 wwl_22_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_5 wbl_21_5 wbl_22_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_5 rwl_22_4 rwl_22_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_5 rbl_21_5 rbl_22_5 rc_unit R0=Rrbl C0=Crbl
xgc_22_6 wwl_22_6 wbl_22_6 rwl_22_6 rbl_22_6 sn_22_6 wos_ros_gc
xrc_wwl_22_6 wwl_22_5 wwl_22_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_6 wbl_21_6 wbl_22_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_6 rwl_22_5 rwl_22_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_6 rbl_21_6 rbl_22_6 rc_unit R0=Rrbl C0=Crbl
xgc_22_7 wwl_22_7 wbl_22_7 rwl_22_7 rbl_22_7 sn_22_7 wos_ros_gc
xrc_wwl_22_7 wwl_22_6 wwl_22_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_7 wbl_21_7 wbl_22_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_7 rwl_22_6 rwl_22_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_7 rbl_21_7 rbl_22_7 rc_unit R0=Rrbl C0=Crbl
xgc_22_8 wwl_22_8 wbl_22_8 rwl_22_8 rbl_22_8 sn_22_8 wos_ros_gc
xrc_wwl_22_8 wwl_22_7 wwl_22_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_8 wbl_21_8 wbl_22_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_8 rwl_22_7 rwl_22_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_8 rbl_21_8 rbl_22_8 rc_unit R0=Rrbl C0=Crbl
xgc_22_9 wwl_22_9 wbl_22_9 rwl_22_9 rbl_22_9 sn_22_9 wos_ros_gc
xrc_wwl_22_9 wwl_22_8 wwl_22_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_9 wbl_21_9 wbl_22_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_9 rwl_22_8 rwl_22_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_9 rbl_21_9 rbl_22_9 rc_unit R0=Rrbl C0=Crbl
xgc_22_10 wwl_22_10 wbl_22_10 rwl_22_10 rbl_22_10 sn_22_10 wos_ros_gc
xrc_wwl_22_10 wwl_22_9 wwl_22_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_10 wbl_21_10 wbl_22_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_10 rwl_22_9 rwl_22_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_10 rbl_21_10 rbl_22_10 rc_unit R0=Rrbl C0=Crbl
xgc_22_11 wwl_22_11 wbl_22_11 rwl_22_11 rbl_22_11 sn_22_11 wos_ros_gc
xrc_wwl_22_11 wwl_22_10 wwl_22_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_11 wbl_21_11 wbl_22_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_11 rwl_22_10 rwl_22_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_11 rbl_21_11 rbl_22_11 rc_unit R0=Rrbl C0=Crbl
xgc_22_12 wwl_22_12 wbl_22_12 rwl_22_12 rbl_22_12 sn_22_12 wos_ros_gc
xrc_wwl_22_12 wwl_22_11 wwl_22_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_12 wbl_21_12 wbl_22_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_12 rwl_22_11 rwl_22_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_12 rbl_21_12 rbl_22_12 rc_unit R0=Rrbl C0=Crbl
xgc_22_13 wwl_22_13 wbl_22_13 rwl_22_13 rbl_22_13 sn_22_13 wos_ros_gc
xrc_wwl_22_13 wwl_22_12 wwl_22_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_13 wbl_21_13 wbl_22_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_13 rwl_22_12 rwl_22_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_13 rbl_21_13 rbl_22_13 rc_unit R0=Rrbl C0=Crbl
xgc_22_14 wwl_22_14 wbl_22_14 rwl_22_14 rbl_22_14 sn_22_14 wos_ros_gc
xrc_wwl_22_14 wwl_22_13 wwl_22_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_14 wbl_21_14 wbl_22_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_14 rwl_22_13 rwl_22_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_14 rbl_21_14 rbl_22_14 rc_unit R0=Rrbl C0=Crbl
xgc_22_15 wwl_22_15 wbl_22_15 rwl_22_15 rbl_22_15 sn_22_15 wos_ros_gc
xrc_wwl_22_15 wwl_22_14 wwl_22_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_15 wbl_21_15 wbl_22_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_15 rwl_22_14 rwl_22_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_15 rbl_21_15 rbl_22_15 rc_unit R0=Rrbl C0=Crbl
xgc_22_16 wwl_22_16 wbl_22_16 rwl_22_16 rbl_22_16 sn_22_16 wos_ros_gc
xrc_wwl_22_16 wwl_22_15 wwl_22_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_16 wbl_21_16 wbl_22_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_16 rwl_22_15 rwl_22_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_16 rbl_21_16 rbl_22_16 rc_unit R0=Rrbl C0=Crbl
xgc_22_17 wwl_22_17 wbl_22_17 rwl_22_17 rbl_22_17 sn_22_17 wos_ros_gc
xrc_wwl_22_17 wwl_22_16 wwl_22_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_17 wbl_21_17 wbl_22_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_17 rwl_22_16 rwl_22_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_17 rbl_21_17 rbl_22_17 rc_unit R0=Rrbl C0=Crbl
xgc_22_18 wwl_22_18 wbl_22_18 rwl_22_18 rbl_22_18 sn_22_18 wos_ros_gc
xrc_wwl_22_18 wwl_22_17 wwl_22_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_18 wbl_21_18 wbl_22_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_18 rwl_22_17 rwl_22_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_18 rbl_21_18 rbl_22_18 rc_unit R0=Rrbl C0=Crbl
xgc_22_19 wwl_22_19 wbl_22_19 rwl_22_19 rbl_22_19 sn_22_19 wos_ros_gc
xrc_wwl_22_19 wwl_22_18 wwl_22_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_19 wbl_21_19 wbl_22_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_19 rwl_22_18 rwl_22_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_19 rbl_21_19 rbl_22_19 rc_unit R0=Rrbl C0=Crbl
xgc_22_20 wwl_22_20 wbl_22_20 rwl_22_20 rbl_22_20 sn_22_20 wos_ros_gc
xrc_wwl_22_20 wwl_22_19 wwl_22_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_20 wbl_21_20 wbl_22_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_20 rwl_22_19 rwl_22_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_20 rbl_21_20 rbl_22_20 rc_unit R0=Rrbl C0=Crbl
xgc_22_21 wwl_22_21 wbl_22_21 rwl_22_21 rbl_22_21 sn_22_21 wos_ros_gc
xrc_wwl_22_21 wwl_22_20 wwl_22_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_21 wbl_21_21 wbl_22_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_21 rwl_22_20 rwl_22_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_21 rbl_21_21 rbl_22_21 rc_unit R0=Rrbl C0=Crbl
xgc_22_22 wwl_22_22 wbl_22_22 rwl_22_22 rbl_22_22 sn_22_22 wos_ros_gc
xrc_wwl_22_22 wwl_22_21 wwl_22_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_22 wbl_21_22 wbl_22_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_22 rwl_22_21 rwl_22_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_22 rbl_21_22 rbl_22_22 rc_unit R0=Rrbl C0=Crbl
xgc_22_23 wwl_22_23 wbl_22_23 rwl_22_23 rbl_22_23 sn_22_23 wos_ros_gc
xrc_wwl_22_23 wwl_22_22 wwl_22_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_23 wbl_21_23 wbl_22_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_23 rwl_22_22 rwl_22_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_23 rbl_21_23 rbl_22_23 rc_unit R0=Rrbl C0=Crbl
xgc_22_24 wwl_22_24 wbl_22_24 rwl_22_24 rbl_22_24 sn_22_24 wos_ros_gc
xrc_wwl_22_24 wwl_22_23 wwl_22_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_24 wbl_21_24 wbl_22_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_24 rwl_22_23 rwl_22_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_24 rbl_21_24 rbl_22_24 rc_unit R0=Rrbl C0=Crbl
xgc_22_25 wwl_22_25 wbl_22_25 rwl_22_25 rbl_22_25 sn_22_25 wos_ros_gc
xrc_wwl_22_25 wwl_22_24 wwl_22_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_25 wbl_21_25 wbl_22_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_25 rwl_22_24 rwl_22_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_25 rbl_21_25 rbl_22_25 rc_unit R0=Rrbl C0=Crbl
xgc_22_26 wwl_22_26 wbl_22_26 rwl_22_26 rbl_22_26 sn_22_26 wos_ros_gc
xrc_wwl_22_26 wwl_22_25 wwl_22_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_26 wbl_21_26 wbl_22_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_26 rwl_22_25 rwl_22_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_26 rbl_21_26 rbl_22_26 rc_unit R0=Rrbl C0=Crbl
xgc_22_27 wwl_22_27 wbl_22_27 rwl_22_27 rbl_22_27 sn_22_27 wos_ros_gc
xrc_wwl_22_27 wwl_22_26 wwl_22_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_27 wbl_21_27 wbl_22_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_27 rwl_22_26 rwl_22_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_27 rbl_21_27 rbl_22_27 rc_unit R0=Rrbl C0=Crbl
xgc_22_28 wwl_22_28 wbl_22_28 rwl_22_28 rbl_22_28 sn_22_28 wos_ros_gc
xrc_wwl_22_28 wwl_22_27 wwl_22_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_28 wbl_21_28 wbl_22_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_28 rwl_22_27 rwl_22_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_28 rbl_21_28 rbl_22_28 rc_unit R0=Rrbl C0=Crbl
xgc_22_29 wwl_22_29 wbl_22_29 rwl_22_29 rbl_22_29 sn_22_29 wos_ros_gc
xrc_wwl_22_29 wwl_22_28 wwl_22_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_29 wbl_21_29 wbl_22_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_29 rwl_22_28 rwl_22_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_29 rbl_21_29 rbl_22_29 rc_unit R0=Rrbl C0=Crbl
xgc_22_30 wwl_22_30 wbl_22_30 rwl_22_30 rbl_22_30 sn_22_30 wos_ros_gc
xrc_wwl_22_30 wwl_22_29 wwl_22_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_30 wbl_21_30 wbl_22_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_30 rwl_22_29 rwl_22_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_30 rbl_21_30 rbl_22_30 rc_unit R0=Rrbl C0=Crbl
xgc_22_31 wwl_22_31 wbl_22_31 rwl_22_31 rbl_22_31 sn_22_31 wos_ros_gc
xrc_wwl_22_31 wwl_22_30 wwl_22_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_22_31 wbl_21_31 wbl_22_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_22_31 rwl_22_30 rwl_22_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_22_31 rbl_21_31 rbl_22_31 rc_unit R0=Rrbl C0=Crbl
xgc_23_0 wwl_23_0 wbl_23_0 rwl_23_0 rbl_23_0 sn_23_0 wos_ros_gc
xrc_wwl_23_0 wwl_23 wwl_23_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_0 wbl_22_0 wbl_23_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_0 rwl_23 rwl_23_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_0 rbl_22_0 rbl_23_0 rc_unit R0=Rrbl C0=Crbl
xgc_23_1 wwl_23_1 wbl_23_1 rwl_23_1 rbl_23_1 sn_23_1 wos_ros_gc
xrc_wwl_23_1 wwl_23_0 wwl_23_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_1 wbl_22_1 wbl_23_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_1 rwl_23_0 rwl_23_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_1 rbl_22_1 rbl_23_1 rc_unit R0=Rrbl C0=Crbl
xgc_23_2 wwl_23_2 wbl_23_2 rwl_23_2 rbl_23_2 sn_23_2 wos_ros_gc
xrc_wwl_23_2 wwl_23_1 wwl_23_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_2 wbl_22_2 wbl_23_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_2 rwl_23_1 rwl_23_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_2 rbl_22_2 rbl_23_2 rc_unit R0=Rrbl C0=Crbl
xgc_23_3 wwl_23_3 wbl_23_3 rwl_23_3 rbl_23_3 sn_23_3 wos_ros_gc
xrc_wwl_23_3 wwl_23_2 wwl_23_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_3 wbl_22_3 wbl_23_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_3 rwl_23_2 rwl_23_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_3 rbl_22_3 rbl_23_3 rc_unit R0=Rrbl C0=Crbl
xgc_23_4 wwl_23_4 wbl_23_4 rwl_23_4 rbl_23_4 sn_23_4 wos_ros_gc
xrc_wwl_23_4 wwl_23_3 wwl_23_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_4 wbl_22_4 wbl_23_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_4 rwl_23_3 rwl_23_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_4 rbl_22_4 rbl_23_4 rc_unit R0=Rrbl C0=Crbl
xgc_23_5 wwl_23_5 wbl_23_5 rwl_23_5 rbl_23_5 sn_23_5 wos_ros_gc
xrc_wwl_23_5 wwl_23_4 wwl_23_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_5 wbl_22_5 wbl_23_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_5 rwl_23_4 rwl_23_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_5 rbl_22_5 rbl_23_5 rc_unit R0=Rrbl C0=Crbl
xgc_23_6 wwl_23_6 wbl_23_6 rwl_23_6 rbl_23_6 sn_23_6 wos_ros_gc
xrc_wwl_23_6 wwl_23_5 wwl_23_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_6 wbl_22_6 wbl_23_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_6 rwl_23_5 rwl_23_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_6 rbl_22_6 rbl_23_6 rc_unit R0=Rrbl C0=Crbl
xgc_23_7 wwl_23_7 wbl_23_7 rwl_23_7 rbl_23_7 sn_23_7 wos_ros_gc
xrc_wwl_23_7 wwl_23_6 wwl_23_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_7 wbl_22_7 wbl_23_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_7 rwl_23_6 rwl_23_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_7 rbl_22_7 rbl_23_7 rc_unit R0=Rrbl C0=Crbl
xgc_23_8 wwl_23_8 wbl_23_8 rwl_23_8 rbl_23_8 sn_23_8 wos_ros_gc
xrc_wwl_23_8 wwl_23_7 wwl_23_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_8 wbl_22_8 wbl_23_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_8 rwl_23_7 rwl_23_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_8 rbl_22_8 rbl_23_8 rc_unit R0=Rrbl C0=Crbl
xgc_23_9 wwl_23_9 wbl_23_9 rwl_23_9 rbl_23_9 sn_23_9 wos_ros_gc
xrc_wwl_23_9 wwl_23_8 wwl_23_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_9 wbl_22_9 wbl_23_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_9 rwl_23_8 rwl_23_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_9 rbl_22_9 rbl_23_9 rc_unit R0=Rrbl C0=Crbl
xgc_23_10 wwl_23_10 wbl_23_10 rwl_23_10 rbl_23_10 sn_23_10 wos_ros_gc
xrc_wwl_23_10 wwl_23_9 wwl_23_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_10 wbl_22_10 wbl_23_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_10 rwl_23_9 rwl_23_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_10 rbl_22_10 rbl_23_10 rc_unit R0=Rrbl C0=Crbl
xgc_23_11 wwl_23_11 wbl_23_11 rwl_23_11 rbl_23_11 sn_23_11 wos_ros_gc
xrc_wwl_23_11 wwl_23_10 wwl_23_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_11 wbl_22_11 wbl_23_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_11 rwl_23_10 rwl_23_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_11 rbl_22_11 rbl_23_11 rc_unit R0=Rrbl C0=Crbl
xgc_23_12 wwl_23_12 wbl_23_12 rwl_23_12 rbl_23_12 sn_23_12 wos_ros_gc
xrc_wwl_23_12 wwl_23_11 wwl_23_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_12 wbl_22_12 wbl_23_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_12 rwl_23_11 rwl_23_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_12 rbl_22_12 rbl_23_12 rc_unit R0=Rrbl C0=Crbl
xgc_23_13 wwl_23_13 wbl_23_13 rwl_23_13 rbl_23_13 sn_23_13 wos_ros_gc
xrc_wwl_23_13 wwl_23_12 wwl_23_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_13 wbl_22_13 wbl_23_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_13 rwl_23_12 rwl_23_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_13 rbl_22_13 rbl_23_13 rc_unit R0=Rrbl C0=Crbl
xgc_23_14 wwl_23_14 wbl_23_14 rwl_23_14 rbl_23_14 sn_23_14 wos_ros_gc
xrc_wwl_23_14 wwl_23_13 wwl_23_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_14 wbl_22_14 wbl_23_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_14 rwl_23_13 rwl_23_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_14 rbl_22_14 rbl_23_14 rc_unit R0=Rrbl C0=Crbl
xgc_23_15 wwl_23_15 wbl_23_15 rwl_23_15 rbl_23_15 sn_23_15 wos_ros_gc
xrc_wwl_23_15 wwl_23_14 wwl_23_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_15 wbl_22_15 wbl_23_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_15 rwl_23_14 rwl_23_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_15 rbl_22_15 rbl_23_15 rc_unit R0=Rrbl C0=Crbl
xgc_23_16 wwl_23_16 wbl_23_16 rwl_23_16 rbl_23_16 sn_23_16 wos_ros_gc
xrc_wwl_23_16 wwl_23_15 wwl_23_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_16 wbl_22_16 wbl_23_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_16 rwl_23_15 rwl_23_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_16 rbl_22_16 rbl_23_16 rc_unit R0=Rrbl C0=Crbl
xgc_23_17 wwl_23_17 wbl_23_17 rwl_23_17 rbl_23_17 sn_23_17 wos_ros_gc
xrc_wwl_23_17 wwl_23_16 wwl_23_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_17 wbl_22_17 wbl_23_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_17 rwl_23_16 rwl_23_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_17 rbl_22_17 rbl_23_17 rc_unit R0=Rrbl C0=Crbl
xgc_23_18 wwl_23_18 wbl_23_18 rwl_23_18 rbl_23_18 sn_23_18 wos_ros_gc
xrc_wwl_23_18 wwl_23_17 wwl_23_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_18 wbl_22_18 wbl_23_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_18 rwl_23_17 rwl_23_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_18 rbl_22_18 rbl_23_18 rc_unit R0=Rrbl C0=Crbl
xgc_23_19 wwl_23_19 wbl_23_19 rwl_23_19 rbl_23_19 sn_23_19 wos_ros_gc
xrc_wwl_23_19 wwl_23_18 wwl_23_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_19 wbl_22_19 wbl_23_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_19 rwl_23_18 rwl_23_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_19 rbl_22_19 rbl_23_19 rc_unit R0=Rrbl C0=Crbl
xgc_23_20 wwl_23_20 wbl_23_20 rwl_23_20 rbl_23_20 sn_23_20 wos_ros_gc
xrc_wwl_23_20 wwl_23_19 wwl_23_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_20 wbl_22_20 wbl_23_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_20 rwl_23_19 rwl_23_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_20 rbl_22_20 rbl_23_20 rc_unit R0=Rrbl C0=Crbl
xgc_23_21 wwl_23_21 wbl_23_21 rwl_23_21 rbl_23_21 sn_23_21 wos_ros_gc
xrc_wwl_23_21 wwl_23_20 wwl_23_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_21 wbl_22_21 wbl_23_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_21 rwl_23_20 rwl_23_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_21 rbl_22_21 rbl_23_21 rc_unit R0=Rrbl C0=Crbl
xgc_23_22 wwl_23_22 wbl_23_22 rwl_23_22 rbl_23_22 sn_23_22 wos_ros_gc
xrc_wwl_23_22 wwl_23_21 wwl_23_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_22 wbl_22_22 wbl_23_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_22 rwl_23_21 rwl_23_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_22 rbl_22_22 rbl_23_22 rc_unit R0=Rrbl C0=Crbl
xgc_23_23 wwl_23_23 wbl_23_23 rwl_23_23 rbl_23_23 sn_23_23 wos_ros_gc
xrc_wwl_23_23 wwl_23_22 wwl_23_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_23 wbl_22_23 wbl_23_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_23 rwl_23_22 rwl_23_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_23 rbl_22_23 rbl_23_23 rc_unit R0=Rrbl C0=Crbl
xgc_23_24 wwl_23_24 wbl_23_24 rwl_23_24 rbl_23_24 sn_23_24 wos_ros_gc
xrc_wwl_23_24 wwl_23_23 wwl_23_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_24 wbl_22_24 wbl_23_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_24 rwl_23_23 rwl_23_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_24 rbl_22_24 rbl_23_24 rc_unit R0=Rrbl C0=Crbl
xgc_23_25 wwl_23_25 wbl_23_25 rwl_23_25 rbl_23_25 sn_23_25 wos_ros_gc
xrc_wwl_23_25 wwl_23_24 wwl_23_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_25 wbl_22_25 wbl_23_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_25 rwl_23_24 rwl_23_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_25 rbl_22_25 rbl_23_25 rc_unit R0=Rrbl C0=Crbl
xgc_23_26 wwl_23_26 wbl_23_26 rwl_23_26 rbl_23_26 sn_23_26 wos_ros_gc
xrc_wwl_23_26 wwl_23_25 wwl_23_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_26 wbl_22_26 wbl_23_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_26 rwl_23_25 rwl_23_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_26 rbl_22_26 rbl_23_26 rc_unit R0=Rrbl C0=Crbl
xgc_23_27 wwl_23_27 wbl_23_27 rwl_23_27 rbl_23_27 sn_23_27 wos_ros_gc
xrc_wwl_23_27 wwl_23_26 wwl_23_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_27 wbl_22_27 wbl_23_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_27 rwl_23_26 rwl_23_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_27 rbl_22_27 rbl_23_27 rc_unit R0=Rrbl C0=Crbl
xgc_23_28 wwl_23_28 wbl_23_28 rwl_23_28 rbl_23_28 sn_23_28 wos_ros_gc
xrc_wwl_23_28 wwl_23_27 wwl_23_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_28 wbl_22_28 wbl_23_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_28 rwl_23_27 rwl_23_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_28 rbl_22_28 rbl_23_28 rc_unit R0=Rrbl C0=Crbl
xgc_23_29 wwl_23_29 wbl_23_29 rwl_23_29 rbl_23_29 sn_23_29 wos_ros_gc
xrc_wwl_23_29 wwl_23_28 wwl_23_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_29 wbl_22_29 wbl_23_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_29 rwl_23_28 rwl_23_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_29 rbl_22_29 rbl_23_29 rc_unit R0=Rrbl C0=Crbl
xgc_23_30 wwl_23_30 wbl_23_30 rwl_23_30 rbl_23_30 sn_23_30 wos_ros_gc
xrc_wwl_23_30 wwl_23_29 wwl_23_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_30 wbl_22_30 wbl_23_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_30 rwl_23_29 rwl_23_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_30 rbl_22_30 rbl_23_30 rc_unit R0=Rrbl C0=Crbl
xgc_23_31 wwl_23_31 wbl_23_31 rwl_23_31 rbl_23_31 sn_23_31 wos_ros_gc
xrc_wwl_23_31 wwl_23_30 wwl_23_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_23_31 wbl_22_31 wbl_23_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_23_31 rwl_23_30 rwl_23_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_23_31 rbl_22_31 rbl_23_31 rc_unit R0=Rrbl C0=Crbl
xgc_24_0 wwl_24_0 wbl_24_0 rwl_24_0 rbl_24_0 sn_24_0 wos_ros_gc
xrc_wwl_24_0 wwl_24 wwl_24_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_0 wbl_23_0 wbl_24_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_0 rwl_24 rwl_24_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_0 rbl_23_0 rbl_24_0 rc_unit R0=Rrbl C0=Crbl
xgc_24_1 wwl_24_1 wbl_24_1 rwl_24_1 rbl_24_1 sn_24_1 wos_ros_gc
xrc_wwl_24_1 wwl_24_0 wwl_24_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_1 wbl_23_1 wbl_24_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_1 rwl_24_0 rwl_24_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_1 rbl_23_1 rbl_24_1 rc_unit R0=Rrbl C0=Crbl
xgc_24_2 wwl_24_2 wbl_24_2 rwl_24_2 rbl_24_2 sn_24_2 wos_ros_gc
xrc_wwl_24_2 wwl_24_1 wwl_24_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_2 wbl_23_2 wbl_24_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_2 rwl_24_1 rwl_24_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_2 rbl_23_2 rbl_24_2 rc_unit R0=Rrbl C0=Crbl
xgc_24_3 wwl_24_3 wbl_24_3 rwl_24_3 rbl_24_3 sn_24_3 wos_ros_gc
xrc_wwl_24_3 wwl_24_2 wwl_24_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_3 wbl_23_3 wbl_24_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_3 rwl_24_2 rwl_24_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_3 rbl_23_3 rbl_24_3 rc_unit R0=Rrbl C0=Crbl
xgc_24_4 wwl_24_4 wbl_24_4 rwl_24_4 rbl_24_4 sn_24_4 wos_ros_gc
xrc_wwl_24_4 wwl_24_3 wwl_24_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_4 wbl_23_4 wbl_24_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_4 rwl_24_3 rwl_24_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_4 rbl_23_4 rbl_24_4 rc_unit R0=Rrbl C0=Crbl
xgc_24_5 wwl_24_5 wbl_24_5 rwl_24_5 rbl_24_5 sn_24_5 wos_ros_gc
xrc_wwl_24_5 wwl_24_4 wwl_24_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_5 wbl_23_5 wbl_24_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_5 rwl_24_4 rwl_24_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_5 rbl_23_5 rbl_24_5 rc_unit R0=Rrbl C0=Crbl
xgc_24_6 wwl_24_6 wbl_24_6 rwl_24_6 rbl_24_6 sn_24_6 wos_ros_gc
xrc_wwl_24_6 wwl_24_5 wwl_24_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_6 wbl_23_6 wbl_24_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_6 rwl_24_5 rwl_24_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_6 rbl_23_6 rbl_24_6 rc_unit R0=Rrbl C0=Crbl
xgc_24_7 wwl_24_7 wbl_24_7 rwl_24_7 rbl_24_7 sn_24_7 wos_ros_gc
xrc_wwl_24_7 wwl_24_6 wwl_24_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_7 wbl_23_7 wbl_24_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_7 rwl_24_6 rwl_24_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_7 rbl_23_7 rbl_24_7 rc_unit R0=Rrbl C0=Crbl
xgc_24_8 wwl_24_8 wbl_24_8 rwl_24_8 rbl_24_8 sn_24_8 wos_ros_gc
xrc_wwl_24_8 wwl_24_7 wwl_24_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_8 wbl_23_8 wbl_24_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_8 rwl_24_7 rwl_24_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_8 rbl_23_8 rbl_24_8 rc_unit R0=Rrbl C0=Crbl
xgc_24_9 wwl_24_9 wbl_24_9 rwl_24_9 rbl_24_9 sn_24_9 wos_ros_gc
xrc_wwl_24_9 wwl_24_8 wwl_24_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_9 wbl_23_9 wbl_24_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_9 rwl_24_8 rwl_24_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_9 rbl_23_9 rbl_24_9 rc_unit R0=Rrbl C0=Crbl
xgc_24_10 wwl_24_10 wbl_24_10 rwl_24_10 rbl_24_10 sn_24_10 wos_ros_gc
xrc_wwl_24_10 wwl_24_9 wwl_24_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_10 wbl_23_10 wbl_24_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_10 rwl_24_9 rwl_24_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_10 rbl_23_10 rbl_24_10 rc_unit R0=Rrbl C0=Crbl
xgc_24_11 wwl_24_11 wbl_24_11 rwl_24_11 rbl_24_11 sn_24_11 wos_ros_gc
xrc_wwl_24_11 wwl_24_10 wwl_24_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_11 wbl_23_11 wbl_24_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_11 rwl_24_10 rwl_24_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_11 rbl_23_11 rbl_24_11 rc_unit R0=Rrbl C0=Crbl
xgc_24_12 wwl_24_12 wbl_24_12 rwl_24_12 rbl_24_12 sn_24_12 wos_ros_gc
xrc_wwl_24_12 wwl_24_11 wwl_24_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_12 wbl_23_12 wbl_24_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_12 rwl_24_11 rwl_24_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_12 rbl_23_12 rbl_24_12 rc_unit R0=Rrbl C0=Crbl
xgc_24_13 wwl_24_13 wbl_24_13 rwl_24_13 rbl_24_13 sn_24_13 wos_ros_gc
xrc_wwl_24_13 wwl_24_12 wwl_24_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_13 wbl_23_13 wbl_24_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_13 rwl_24_12 rwl_24_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_13 rbl_23_13 rbl_24_13 rc_unit R0=Rrbl C0=Crbl
xgc_24_14 wwl_24_14 wbl_24_14 rwl_24_14 rbl_24_14 sn_24_14 wos_ros_gc
xrc_wwl_24_14 wwl_24_13 wwl_24_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_14 wbl_23_14 wbl_24_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_14 rwl_24_13 rwl_24_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_14 rbl_23_14 rbl_24_14 rc_unit R0=Rrbl C0=Crbl
xgc_24_15 wwl_24_15 wbl_24_15 rwl_24_15 rbl_24_15 sn_24_15 wos_ros_gc
xrc_wwl_24_15 wwl_24_14 wwl_24_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_15 wbl_23_15 wbl_24_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_15 rwl_24_14 rwl_24_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_15 rbl_23_15 rbl_24_15 rc_unit R0=Rrbl C0=Crbl
xgc_24_16 wwl_24_16 wbl_24_16 rwl_24_16 rbl_24_16 sn_24_16 wos_ros_gc
xrc_wwl_24_16 wwl_24_15 wwl_24_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_16 wbl_23_16 wbl_24_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_16 rwl_24_15 rwl_24_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_16 rbl_23_16 rbl_24_16 rc_unit R0=Rrbl C0=Crbl
xgc_24_17 wwl_24_17 wbl_24_17 rwl_24_17 rbl_24_17 sn_24_17 wos_ros_gc
xrc_wwl_24_17 wwl_24_16 wwl_24_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_17 wbl_23_17 wbl_24_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_17 rwl_24_16 rwl_24_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_17 rbl_23_17 rbl_24_17 rc_unit R0=Rrbl C0=Crbl
xgc_24_18 wwl_24_18 wbl_24_18 rwl_24_18 rbl_24_18 sn_24_18 wos_ros_gc
xrc_wwl_24_18 wwl_24_17 wwl_24_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_18 wbl_23_18 wbl_24_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_18 rwl_24_17 rwl_24_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_18 rbl_23_18 rbl_24_18 rc_unit R0=Rrbl C0=Crbl
xgc_24_19 wwl_24_19 wbl_24_19 rwl_24_19 rbl_24_19 sn_24_19 wos_ros_gc
xrc_wwl_24_19 wwl_24_18 wwl_24_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_19 wbl_23_19 wbl_24_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_19 rwl_24_18 rwl_24_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_19 rbl_23_19 rbl_24_19 rc_unit R0=Rrbl C0=Crbl
xgc_24_20 wwl_24_20 wbl_24_20 rwl_24_20 rbl_24_20 sn_24_20 wos_ros_gc
xrc_wwl_24_20 wwl_24_19 wwl_24_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_20 wbl_23_20 wbl_24_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_20 rwl_24_19 rwl_24_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_20 rbl_23_20 rbl_24_20 rc_unit R0=Rrbl C0=Crbl
xgc_24_21 wwl_24_21 wbl_24_21 rwl_24_21 rbl_24_21 sn_24_21 wos_ros_gc
xrc_wwl_24_21 wwl_24_20 wwl_24_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_21 wbl_23_21 wbl_24_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_21 rwl_24_20 rwl_24_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_21 rbl_23_21 rbl_24_21 rc_unit R0=Rrbl C0=Crbl
xgc_24_22 wwl_24_22 wbl_24_22 rwl_24_22 rbl_24_22 sn_24_22 wos_ros_gc
xrc_wwl_24_22 wwl_24_21 wwl_24_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_22 wbl_23_22 wbl_24_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_22 rwl_24_21 rwl_24_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_22 rbl_23_22 rbl_24_22 rc_unit R0=Rrbl C0=Crbl
xgc_24_23 wwl_24_23 wbl_24_23 rwl_24_23 rbl_24_23 sn_24_23 wos_ros_gc
xrc_wwl_24_23 wwl_24_22 wwl_24_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_23 wbl_23_23 wbl_24_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_23 rwl_24_22 rwl_24_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_23 rbl_23_23 rbl_24_23 rc_unit R0=Rrbl C0=Crbl
xgc_24_24 wwl_24_24 wbl_24_24 rwl_24_24 rbl_24_24 sn_24_24 wos_ros_gc
xrc_wwl_24_24 wwl_24_23 wwl_24_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_24 wbl_23_24 wbl_24_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_24 rwl_24_23 rwl_24_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_24 rbl_23_24 rbl_24_24 rc_unit R0=Rrbl C0=Crbl
xgc_24_25 wwl_24_25 wbl_24_25 rwl_24_25 rbl_24_25 sn_24_25 wos_ros_gc
xrc_wwl_24_25 wwl_24_24 wwl_24_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_25 wbl_23_25 wbl_24_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_25 rwl_24_24 rwl_24_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_25 rbl_23_25 rbl_24_25 rc_unit R0=Rrbl C0=Crbl
xgc_24_26 wwl_24_26 wbl_24_26 rwl_24_26 rbl_24_26 sn_24_26 wos_ros_gc
xrc_wwl_24_26 wwl_24_25 wwl_24_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_26 wbl_23_26 wbl_24_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_26 rwl_24_25 rwl_24_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_26 rbl_23_26 rbl_24_26 rc_unit R0=Rrbl C0=Crbl
xgc_24_27 wwl_24_27 wbl_24_27 rwl_24_27 rbl_24_27 sn_24_27 wos_ros_gc
xrc_wwl_24_27 wwl_24_26 wwl_24_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_27 wbl_23_27 wbl_24_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_27 rwl_24_26 rwl_24_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_27 rbl_23_27 rbl_24_27 rc_unit R0=Rrbl C0=Crbl
xgc_24_28 wwl_24_28 wbl_24_28 rwl_24_28 rbl_24_28 sn_24_28 wos_ros_gc
xrc_wwl_24_28 wwl_24_27 wwl_24_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_28 wbl_23_28 wbl_24_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_28 rwl_24_27 rwl_24_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_28 rbl_23_28 rbl_24_28 rc_unit R0=Rrbl C0=Crbl
xgc_24_29 wwl_24_29 wbl_24_29 rwl_24_29 rbl_24_29 sn_24_29 wos_ros_gc
xrc_wwl_24_29 wwl_24_28 wwl_24_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_29 wbl_23_29 wbl_24_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_29 rwl_24_28 rwl_24_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_29 rbl_23_29 rbl_24_29 rc_unit R0=Rrbl C0=Crbl
xgc_24_30 wwl_24_30 wbl_24_30 rwl_24_30 rbl_24_30 sn_24_30 wos_ros_gc
xrc_wwl_24_30 wwl_24_29 wwl_24_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_30 wbl_23_30 wbl_24_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_30 rwl_24_29 rwl_24_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_30 rbl_23_30 rbl_24_30 rc_unit R0=Rrbl C0=Crbl
xgc_24_31 wwl_24_31 wbl_24_31 rwl_24_31 rbl_24_31 sn_24_31 wos_ros_gc
xrc_wwl_24_31 wwl_24_30 wwl_24_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_24_31 wbl_23_31 wbl_24_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_24_31 rwl_24_30 rwl_24_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_24_31 rbl_23_31 rbl_24_31 rc_unit R0=Rrbl C0=Crbl
xgc_25_0 wwl_25_0 wbl_25_0 rwl_25_0 rbl_25_0 sn_25_0 wos_ros_gc
xrc_wwl_25_0 wwl_25 wwl_25_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_0 wbl_24_0 wbl_25_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_0 rwl_25 rwl_25_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_0 rbl_24_0 rbl_25_0 rc_unit R0=Rrbl C0=Crbl
xgc_25_1 wwl_25_1 wbl_25_1 rwl_25_1 rbl_25_1 sn_25_1 wos_ros_gc
xrc_wwl_25_1 wwl_25_0 wwl_25_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_1 wbl_24_1 wbl_25_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_1 rwl_25_0 rwl_25_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_1 rbl_24_1 rbl_25_1 rc_unit R0=Rrbl C0=Crbl
xgc_25_2 wwl_25_2 wbl_25_2 rwl_25_2 rbl_25_2 sn_25_2 wos_ros_gc
xrc_wwl_25_2 wwl_25_1 wwl_25_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_2 wbl_24_2 wbl_25_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_2 rwl_25_1 rwl_25_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_2 rbl_24_2 rbl_25_2 rc_unit R0=Rrbl C0=Crbl
xgc_25_3 wwl_25_3 wbl_25_3 rwl_25_3 rbl_25_3 sn_25_3 wos_ros_gc
xrc_wwl_25_3 wwl_25_2 wwl_25_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_3 wbl_24_3 wbl_25_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_3 rwl_25_2 rwl_25_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_3 rbl_24_3 rbl_25_3 rc_unit R0=Rrbl C0=Crbl
xgc_25_4 wwl_25_4 wbl_25_4 rwl_25_4 rbl_25_4 sn_25_4 wos_ros_gc
xrc_wwl_25_4 wwl_25_3 wwl_25_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_4 wbl_24_4 wbl_25_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_4 rwl_25_3 rwl_25_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_4 rbl_24_4 rbl_25_4 rc_unit R0=Rrbl C0=Crbl
xgc_25_5 wwl_25_5 wbl_25_5 rwl_25_5 rbl_25_5 sn_25_5 wos_ros_gc
xrc_wwl_25_5 wwl_25_4 wwl_25_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_5 wbl_24_5 wbl_25_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_5 rwl_25_4 rwl_25_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_5 rbl_24_5 rbl_25_5 rc_unit R0=Rrbl C0=Crbl
xgc_25_6 wwl_25_6 wbl_25_6 rwl_25_6 rbl_25_6 sn_25_6 wos_ros_gc
xrc_wwl_25_6 wwl_25_5 wwl_25_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_6 wbl_24_6 wbl_25_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_6 rwl_25_5 rwl_25_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_6 rbl_24_6 rbl_25_6 rc_unit R0=Rrbl C0=Crbl
xgc_25_7 wwl_25_7 wbl_25_7 rwl_25_7 rbl_25_7 sn_25_7 wos_ros_gc
xrc_wwl_25_7 wwl_25_6 wwl_25_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_7 wbl_24_7 wbl_25_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_7 rwl_25_6 rwl_25_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_7 rbl_24_7 rbl_25_7 rc_unit R0=Rrbl C0=Crbl
xgc_25_8 wwl_25_8 wbl_25_8 rwl_25_8 rbl_25_8 sn_25_8 wos_ros_gc
xrc_wwl_25_8 wwl_25_7 wwl_25_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_8 wbl_24_8 wbl_25_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_8 rwl_25_7 rwl_25_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_8 rbl_24_8 rbl_25_8 rc_unit R0=Rrbl C0=Crbl
xgc_25_9 wwl_25_9 wbl_25_9 rwl_25_9 rbl_25_9 sn_25_9 wos_ros_gc
xrc_wwl_25_9 wwl_25_8 wwl_25_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_9 wbl_24_9 wbl_25_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_9 rwl_25_8 rwl_25_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_9 rbl_24_9 rbl_25_9 rc_unit R0=Rrbl C0=Crbl
xgc_25_10 wwl_25_10 wbl_25_10 rwl_25_10 rbl_25_10 sn_25_10 wos_ros_gc
xrc_wwl_25_10 wwl_25_9 wwl_25_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_10 wbl_24_10 wbl_25_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_10 rwl_25_9 rwl_25_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_10 rbl_24_10 rbl_25_10 rc_unit R0=Rrbl C0=Crbl
xgc_25_11 wwl_25_11 wbl_25_11 rwl_25_11 rbl_25_11 sn_25_11 wos_ros_gc
xrc_wwl_25_11 wwl_25_10 wwl_25_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_11 wbl_24_11 wbl_25_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_11 rwl_25_10 rwl_25_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_11 rbl_24_11 rbl_25_11 rc_unit R0=Rrbl C0=Crbl
xgc_25_12 wwl_25_12 wbl_25_12 rwl_25_12 rbl_25_12 sn_25_12 wos_ros_gc
xrc_wwl_25_12 wwl_25_11 wwl_25_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_12 wbl_24_12 wbl_25_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_12 rwl_25_11 rwl_25_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_12 rbl_24_12 rbl_25_12 rc_unit R0=Rrbl C0=Crbl
xgc_25_13 wwl_25_13 wbl_25_13 rwl_25_13 rbl_25_13 sn_25_13 wos_ros_gc
xrc_wwl_25_13 wwl_25_12 wwl_25_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_13 wbl_24_13 wbl_25_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_13 rwl_25_12 rwl_25_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_13 rbl_24_13 rbl_25_13 rc_unit R0=Rrbl C0=Crbl
xgc_25_14 wwl_25_14 wbl_25_14 rwl_25_14 rbl_25_14 sn_25_14 wos_ros_gc
xrc_wwl_25_14 wwl_25_13 wwl_25_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_14 wbl_24_14 wbl_25_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_14 rwl_25_13 rwl_25_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_14 rbl_24_14 rbl_25_14 rc_unit R0=Rrbl C0=Crbl
xgc_25_15 wwl_25_15 wbl_25_15 rwl_25_15 rbl_25_15 sn_25_15 wos_ros_gc
xrc_wwl_25_15 wwl_25_14 wwl_25_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_15 wbl_24_15 wbl_25_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_15 rwl_25_14 rwl_25_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_15 rbl_24_15 rbl_25_15 rc_unit R0=Rrbl C0=Crbl
xgc_25_16 wwl_25_16 wbl_25_16 rwl_25_16 rbl_25_16 sn_25_16 wos_ros_gc
xrc_wwl_25_16 wwl_25_15 wwl_25_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_16 wbl_24_16 wbl_25_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_16 rwl_25_15 rwl_25_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_16 rbl_24_16 rbl_25_16 rc_unit R0=Rrbl C0=Crbl
xgc_25_17 wwl_25_17 wbl_25_17 rwl_25_17 rbl_25_17 sn_25_17 wos_ros_gc
xrc_wwl_25_17 wwl_25_16 wwl_25_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_17 wbl_24_17 wbl_25_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_17 rwl_25_16 rwl_25_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_17 rbl_24_17 rbl_25_17 rc_unit R0=Rrbl C0=Crbl
xgc_25_18 wwl_25_18 wbl_25_18 rwl_25_18 rbl_25_18 sn_25_18 wos_ros_gc
xrc_wwl_25_18 wwl_25_17 wwl_25_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_18 wbl_24_18 wbl_25_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_18 rwl_25_17 rwl_25_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_18 rbl_24_18 rbl_25_18 rc_unit R0=Rrbl C0=Crbl
xgc_25_19 wwl_25_19 wbl_25_19 rwl_25_19 rbl_25_19 sn_25_19 wos_ros_gc
xrc_wwl_25_19 wwl_25_18 wwl_25_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_19 wbl_24_19 wbl_25_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_19 rwl_25_18 rwl_25_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_19 rbl_24_19 rbl_25_19 rc_unit R0=Rrbl C0=Crbl
xgc_25_20 wwl_25_20 wbl_25_20 rwl_25_20 rbl_25_20 sn_25_20 wos_ros_gc
xrc_wwl_25_20 wwl_25_19 wwl_25_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_20 wbl_24_20 wbl_25_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_20 rwl_25_19 rwl_25_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_20 rbl_24_20 rbl_25_20 rc_unit R0=Rrbl C0=Crbl
xgc_25_21 wwl_25_21 wbl_25_21 rwl_25_21 rbl_25_21 sn_25_21 wos_ros_gc
xrc_wwl_25_21 wwl_25_20 wwl_25_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_21 wbl_24_21 wbl_25_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_21 rwl_25_20 rwl_25_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_21 rbl_24_21 rbl_25_21 rc_unit R0=Rrbl C0=Crbl
xgc_25_22 wwl_25_22 wbl_25_22 rwl_25_22 rbl_25_22 sn_25_22 wos_ros_gc
xrc_wwl_25_22 wwl_25_21 wwl_25_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_22 wbl_24_22 wbl_25_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_22 rwl_25_21 rwl_25_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_22 rbl_24_22 rbl_25_22 rc_unit R0=Rrbl C0=Crbl
xgc_25_23 wwl_25_23 wbl_25_23 rwl_25_23 rbl_25_23 sn_25_23 wos_ros_gc
xrc_wwl_25_23 wwl_25_22 wwl_25_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_23 wbl_24_23 wbl_25_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_23 rwl_25_22 rwl_25_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_23 rbl_24_23 rbl_25_23 rc_unit R0=Rrbl C0=Crbl
xgc_25_24 wwl_25_24 wbl_25_24 rwl_25_24 rbl_25_24 sn_25_24 wos_ros_gc
xrc_wwl_25_24 wwl_25_23 wwl_25_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_24 wbl_24_24 wbl_25_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_24 rwl_25_23 rwl_25_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_24 rbl_24_24 rbl_25_24 rc_unit R0=Rrbl C0=Crbl
xgc_25_25 wwl_25_25 wbl_25_25 rwl_25_25 rbl_25_25 sn_25_25 wos_ros_gc
xrc_wwl_25_25 wwl_25_24 wwl_25_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_25 wbl_24_25 wbl_25_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_25 rwl_25_24 rwl_25_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_25 rbl_24_25 rbl_25_25 rc_unit R0=Rrbl C0=Crbl
xgc_25_26 wwl_25_26 wbl_25_26 rwl_25_26 rbl_25_26 sn_25_26 wos_ros_gc
xrc_wwl_25_26 wwl_25_25 wwl_25_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_26 wbl_24_26 wbl_25_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_26 rwl_25_25 rwl_25_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_26 rbl_24_26 rbl_25_26 rc_unit R0=Rrbl C0=Crbl
xgc_25_27 wwl_25_27 wbl_25_27 rwl_25_27 rbl_25_27 sn_25_27 wos_ros_gc
xrc_wwl_25_27 wwl_25_26 wwl_25_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_27 wbl_24_27 wbl_25_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_27 rwl_25_26 rwl_25_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_27 rbl_24_27 rbl_25_27 rc_unit R0=Rrbl C0=Crbl
xgc_25_28 wwl_25_28 wbl_25_28 rwl_25_28 rbl_25_28 sn_25_28 wos_ros_gc
xrc_wwl_25_28 wwl_25_27 wwl_25_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_28 wbl_24_28 wbl_25_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_28 rwl_25_27 rwl_25_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_28 rbl_24_28 rbl_25_28 rc_unit R0=Rrbl C0=Crbl
xgc_25_29 wwl_25_29 wbl_25_29 rwl_25_29 rbl_25_29 sn_25_29 wos_ros_gc
xrc_wwl_25_29 wwl_25_28 wwl_25_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_29 wbl_24_29 wbl_25_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_29 rwl_25_28 rwl_25_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_29 rbl_24_29 rbl_25_29 rc_unit R0=Rrbl C0=Crbl
xgc_25_30 wwl_25_30 wbl_25_30 rwl_25_30 rbl_25_30 sn_25_30 wos_ros_gc
xrc_wwl_25_30 wwl_25_29 wwl_25_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_30 wbl_24_30 wbl_25_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_30 rwl_25_29 rwl_25_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_30 rbl_24_30 rbl_25_30 rc_unit R0=Rrbl C0=Crbl
xgc_25_31 wwl_25_31 wbl_25_31 rwl_25_31 rbl_25_31 sn_25_31 wos_ros_gc
xrc_wwl_25_31 wwl_25_30 wwl_25_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_25_31 wbl_24_31 wbl_25_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_25_31 rwl_25_30 rwl_25_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_25_31 rbl_24_31 rbl_25_31 rc_unit R0=Rrbl C0=Crbl
xgc_26_0 wwl_26_0 wbl_26_0 rwl_26_0 rbl_26_0 sn_26_0 wos_ros_gc
xrc_wwl_26_0 wwl_26 wwl_26_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_0 wbl_25_0 wbl_26_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_0 rwl_26 rwl_26_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_0 rbl_25_0 rbl_26_0 rc_unit R0=Rrbl C0=Crbl
xgc_26_1 wwl_26_1 wbl_26_1 rwl_26_1 rbl_26_1 sn_26_1 wos_ros_gc
xrc_wwl_26_1 wwl_26_0 wwl_26_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_1 wbl_25_1 wbl_26_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_1 rwl_26_0 rwl_26_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_1 rbl_25_1 rbl_26_1 rc_unit R0=Rrbl C0=Crbl
xgc_26_2 wwl_26_2 wbl_26_2 rwl_26_2 rbl_26_2 sn_26_2 wos_ros_gc
xrc_wwl_26_2 wwl_26_1 wwl_26_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_2 wbl_25_2 wbl_26_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_2 rwl_26_1 rwl_26_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_2 rbl_25_2 rbl_26_2 rc_unit R0=Rrbl C0=Crbl
xgc_26_3 wwl_26_3 wbl_26_3 rwl_26_3 rbl_26_3 sn_26_3 wos_ros_gc
xrc_wwl_26_3 wwl_26_2 wwl_26_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_3 wbl_25_3 wbl_26_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_3 rwl_26_2 rwl_26_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_3 rbl_25_3 rbl_26_3 rc_unit R0=Rrbl C0=Crbl
xgc_26_4 wwl_26_4 wbl_26_4 rwl_26_4 rbl_26_4 sn_26_4 wos_ros_gc
xrc_wwl_26_4 wwl_26_3 wwl_26_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_4 wbl_25_4 wbl_26_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_4 rwl_26_3 rwl_26_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_4 rbl_25_4 rbl_26_4 rc_unit R0=Rrbl C0=Crbl
xgc_26_5 wwl_26_5 wbl_26_5 rwl_26_5 rbl_26_5 sn_26_5 wos_ros_gc
xrc_wwl_26_5 wwl_26_4 wwl_26_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_5 wbl_25_5 wbl_26_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_5 rwl_26_4 rwl_26_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_5 rbl_25_5 rbl_26_5 rc_unit R0=Rrbl C0=Crbl
xgc_26_6 wwl_26_6 wbl_26_6 rwl_26_6 rbl_26_6 sn_26_6 wos_ros_gc
xrc_wwl_26_6 wwl_26_5 wwl_26_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_6 wbl_25_6 wbl_26_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_6 rwl_26_5 rwl_26_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_6 rbl_25_6 rbl_26_6 rc_unit R0=Rrbl C0=Crbl
xgc_26_7 wwl_26_7 wbl_26_7 rwl_26_7 rbl_26_7 sn_26_7 wos_ros_gc
xrc_wwl_26_7 wwl_26_6 wwl_26_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_7 wbl_25_7 wbl_26_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_7 rwl_26_6 rwl_26_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_7 rbl_25_7 rbl_26_7 rc_unit R0=Rrbl C0=Crbl
xgc_26_8 wwl_26_8 wbl_26_8 rwl_26_8 rbl_26_8 sn_26_8 wos_ros_gc
xrc_wwl_26_8 wwl_26_7 wwl_26_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_8 wbl_25_8 wbl_26_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_8 rwl_26_7 rwl_26_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_8 rbl_25_8 rbl_26_8 rc_unit R0=Rrbl C0=Crbl
xgc_26_9 wwl_26_9 wbl_26_9 rwl_26_9 rbl_26_9 sn_26_9 wos_ros_gc
xrc_wwl_26_9 wwl_26_8 wwl_26_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_9 wbl_25_9 wbl_26_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_9 rwl_26_8 rwl_26_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_9 rbl_25_9 rbl_26_9 rc_unit R0=Rrbl C0=Crbl
xgc_26_10 wwl_26_10 wbl_26_10 rwl_26_10 rbl_26_10 sn_26_10 wos_ros_gc
xrc_wwl_26_10 wwl_26_9 wwl_26_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_10 wbl_25_10 wbl_26_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_10 rwl_26_9 rwl_26_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_10 rbl_25_10 rbl_26_10 rc_unit R0=Rrbl C0=Crbl
xgc_26_11 wwl_26_11 wbl_26_11 rwl_26_11 rbl_26_11 sn_26_11 wos_ros_gc
xrc_wwl_26_11 wwl_26_10 wwl_26_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_11 wbl_25_11 wbl_26_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_11 rwl_26_10 rwl_26_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_11 rbl_25_11 rbl_26_11 rc_unit R0=Rrbl C0=Crbl
xgc_26_12 wwl_26_12 wbl_26_12 rwl_26_12 rbl_26_12 sn_26_12 wos_ros_gc
xrc_wwl_26_12 wwl_26_11 wwl_26_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_12 wbl_25_12 wbl_26_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_12 rwl_26_11 rwl_26_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_12 rbl_25_12 rbl_26_12 rc_unit R0=Rrbl C0=Crbl
xgc_26_13 wwl_26_13 wbl_26_13 rwl_26_13 rbl_26_13 sn_26_13 wos_ros_gc
xrc_wwl_26_13 wwl_26_12 wwl_26_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_13 wbl_25_13 wbl_26_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_13 rwl_26_12 rwl_26_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_13 rbl_25_13 rbl_26_13 rc_unit R0=Rrbl C0=Crbl
xgc_26_14 wwl_26_14 wbl_26_14 rwl_26_14 rbl_26_14 sn_26_14 wos_ros_gc
xrc_wwl_26_14 wwl_26_13 wwl_26_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_14 wbl_25_14 wbl_26_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_14 rwl_26_13 rwl_26_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_14 rbl_25_14 rbl_26_14 rc_unit R0=Rrbl C0=Crbl
xgc_26_15 wwl_26_15 wbl_26_15 rwl_26_15 rbl_26_15 sn_26_15 wos_ros_gc
xrc_wwl_26_15 wwl_26_14 wwl_26_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_15 wbl_25_15 wbl_26_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_15 rwl_26_14 rwl_26_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_15 rbl_25_15 rbl_26_15 rc_unit R0=Rrbl C0=Crbl
xgc_26_16 wwl_26_16 wbl_26_16 rwl_26_16 rbl_26_16 sn_26_16 wos_ros_gc
xrc_wwl_26_16 wwl_26_15 wwl_26_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_16 wbl_25_16 wbl_26_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_16 rwl_26_15 rwl_26_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_16 rbl_25_16 rbl_26_16 rc_unit R0=Rrbl C0=Crbl
xgc_26_17 wwl_26_17 wbl_26_17 rwl_26_17 rbl_26_17 sn_26_17 wos_ros_gc
xrc_wwl_26_17 wwl_26_16 wwl_26_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_17 wbl_25_17 wbl_26_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_17 rwl_26_16 rwl_26_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_17 rbl_25_17 rbl_26_17 rc_unit R0=Rrbl C0=Crbl
xgc_26_18 wwl_26_18 wbl_26_18 rwl_26_18 rbl_26_18 sn_26_18 wos_ros_gc
xrc_wwl_26_18 wwl_26_17 wwl_26_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_18 wbl_25_18 wbl_26_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_18 rwl_26_17 rwl_26_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_18 rbl_25_18 rbl_26_18 rc_unit R0=Rrbl C0=Crbl
xgc_26_19 wwl_26_19 wbl_26_19 rwl_26_19 rbl_26_19 sn_26_19 wos_ros_gc
xrc_wwl_26_19 wwl_26_18 wwl_26_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_19 wbl_25_19 wbl_26_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_19 rwl_26_18 rwl_26_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_19 rbl_25_19 rbl_26_19 rc_unit R0=Rrbl C0=Crbl
xgc_26_20 wwl_26_20 wbl_26_20 rwl_26_20 rbl_26_20 sn_26_20 wos_ros_gc
xrc_wwl_26_20 wwl_26_19 wwl_26_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_20 wbl_25_20 wbl_26_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_20 rwl_26_19 rwl_26_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_20 rbl_25_20 rbl_26_20 rc_unit R0=Rrbl C0=Crbl
xgc_26_21 wwl_26_21 wbl_26_21 rwl_26_21 rbl_26_21 sn_26_21 wos_ros_gc
xrc_wwl_26_21 wwl_26_20 wwl_26_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_21 wbl_25_21 wbl_26_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_21 rwl_26_20 rwl_26_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_21 rbl_25_21 rbl_26_21 rc_unit R0=Rrbl C0=Crbl
xgc_26_22 wwl_26_22 wbl_26_22 rwl_26_22 rbl_26_22 sn_26_22 wos_ros_gc
xrc_wwl_26_22 wwl_26_21 wwl_26_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_22 wbl_25_22 wbl_26_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_22 rwl_26_21 rwl_26_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_22 rbl_25_22 rbl_26_22 rc_unit R0=Rrbl C0=Crbl
xgc_26_23 wwl_26_23 wbl_26_23 rwl_26_23 rbl_26_23 sn_26_23 wos_ros_gc
xrc_wwl_26_23 wwl_26_22 wwl_26_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_23 wbl_25_23 wbl_26_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_23 rwl_26_22 rwl_26_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_23 rbl_25_23 rbl_26_23 rc_unit R0=Rrbl C0=Crbl
xgc_26_24 wwl_26_24 wbl_26_24 rwl_26_24 rbl_26_24 sn_26_24 wos_ros_gc
xrc_wwl_26_24 wwl_26_23 wwl_26_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_24 wbl_25_24 wbl_26_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_24 rwl_26_23 rwl_26_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_24 rbl_25_24 rbl_26_24 rc_unit R0=Rrbl C0=Crbl
xgc_26_25 wwl_26_25 wbl_26_25 rwl_26_25 rbl_26_25 sn_26_25 wos_ros_gc
xrc_wwl_26_25 wwl_26_24 wwl_26_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_25 wbl_25_25 wbl_26_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_25 rwl_26_24 rwl_26_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_25 rbl_25_25 rbl_26_25 rc_unit R0=Rrbl C0=Crbl
xgc_26_26 wwl_26_26 wbl_26_26 rwl_26_26 rbl_26_26 sn_26_26 wos_ros_gc
xrc_wwl_26_26 wwl_26_25 wwl_26_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_26 wbl_25_26 wbl_26_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_26 rwl_26_25 rwl_26_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_26 rbl_25_26 rbl_26_26 rc_unit R0=Rrbl C0=Crbl
xgc_26_27 wwl_26_27 wbl_26_27 rwl_26_27 rbl_26_27 sn_26_27 wos_ros_gc
xrc_wwl_26_27 wwl_26_26 wwl_26_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_27 wbl_25_27 wbl_26_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_27 rwl_26_26 rwl_26_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_27 rbl_25_27 rbl_26_27 rc_unit R0=Rrbl C0=Crbl
xgc_26_28 wwl_26_28 wbl_26_28 rwl_26_28 rbl_26_28 sn_26_28 wos_ros_gc
xrc_wwl_26_28 wwl_26_27 wwl_26_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_28 wbl_25_28 wbl_26_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_28 rwl_26_27 rwl_26_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_28 rbl_25_28 rbl_26_28 rc_unit R0=Rrbl C0=Crbl
xgc_26_29 wwl_26_29 wbl_26_29 rwl_26_29 rbl_26_29 sn_26_29 wos_ros_gc
xrc_wwl_26_29 wwl_26_28 wwl_26_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_29 wbl_25_29 wbl_26_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_29 rwl_26_28 rwl_26_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_29 rbl_25_29 rbl_26_29 rc_unit R0=Rrbl C0=Crbl
xgc_26_30 wwl_26_30 wbl_26_30 rwl_26_30 rbl_26_30 sn_26_30 wos_ros_gc
xrc_wwl_26_30 wwl_26_29 wwl_26_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_30 wbl_25_30 wbl_26_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_30 rwl_26_29 rwl_26_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_30 rbl_25_30 rbl_26_30 rc_unit R0=Rrbl C0=Crbl
xgc_26_31 wwl_26_31 wbl_26_31 rwl_26_31 rbl_26_31 sn_26_31 wos_ros_gc
xrc_wwl_26_31 wwl_26_30 wwl_26_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_26_31 wbl_25_31 wbl_26_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_26_31 rwl_26_30 rwl_26_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_26_31 rbl_25_31 rbl_26_31 rc_unit R0=Rrbl C0=Crbl
xgc_27_0 wwl_27_0 wbl_27_0 rwl_27_0 rbl_27_0 sn_27_0 wos_ros_gc
xrc_wwl_27_0 wwl_27 wwl_27_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_0 wbl_26_0 wbl_27_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_0 rwl_27 rwl_27_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_0 rbl_26_0 rbl_27_0 rc_unit R0=Rrbl C0=Crbl
xgc_27_1 wwl_27_1 wbl_27_1 rwl_27_1 rbl_27_1 sn_27_1 wos_ros_gc
xrc_wwl_27_1 wwl_27_0 wwl_27_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_1 wbl_26_1 wbl_27_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_1 rwl_27_0 rwl_27_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_1 rbl_26_1 rbl_27_1 rc_unit R0=Rrbl C0=Crbl
xgc_27_2 wwl_27_2 wbl_27_2 rwl_27_2 rbl_27_2 sn_27_2 wos_ros_gc
xrc_wwl_27_2 wwl_27_1 wwl_27_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_2 wbl_26_2 wbl_27_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_2 rwl_27_1 rwl_27_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_2 rbl_26_2 rbl_27_2 rc_unit R0=Rrbl C0=Crbl
xgc_27_3 wwl_27_3 wbl_27_3 rwl_27_3 rbl_27_3 sn_27_3 wos_ros_gc
xrc_wwl_27_3 wwl_27_2 wwl_27_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_3 wbl_26_3 wbl_27_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_3 rwl_27_2 rwl_27_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_3 rbl_26_3 rbl_27_3 rc_unit R0=Rrbl C0=Crbl
xgc_27_4 wwl_27_4 wbl_27_4 rwl_27_4 rbl_27_4 sn_27_4 wos_ros_gc
xrc_wwl_27_4 wwl_27_3 wwl_27_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_4 wbl_26_4 wbl_27_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_4 rwl_27_3 rwl_27_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_4 rbl_26_4 rbl_27_4 rc_unit R0=Rrbl C0=Crbl
xgc_27_5 wwl_27_5 wbl_27_5 rwl_27_5 rbl_27_5 sn_27_5 wos_ros_gc
xrc_wwl_27_5 wwl_27_4 wwl_27_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_5 wbl_26_5 wbl_27_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_5 rwl_27_4 rwl_27_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_5 rbl_26_5 rbl_27_5 rc_unit R0=Rrbl C0=Crbl
xgc_27_6 wwl_27_6 wbl_27_6 rwl_27_6 rbl_27_6 sn_27_6 wos_ros_gc
xrc_wwl_27_6 wwl_27_5 wwl_27_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_6 wbl_26_6 wbl_27_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_6 rwl_27_5 rwl_27_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_6 rbl_26_6 rbl_27_6 rc_unit R0=Rrbl C0=Crbl
xgc_27_7 wwl_27_7 wbl_27_7 rwl_27_7 rbl_27_7 sn_27_7 wos_ros_gc
xrc_wwl_27_7 wwl_27_6 wwl_27_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_7 wbl_26_7 wbl_27_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_7 rwl_27_6 rwl_27_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_7 rbl_26_7 rbl_27_7 rc_unit R0=Rrbl C0=Crbl
xgc_27_8 wwl_27_8 wbl_27_8 rwl_27_8 rbl_27_8 sn_27_8 wos_ros_gc
xrc_wwl_27_8 wwl_27_7 wwl_27_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_8 wbl_26_8 wbl_27_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_8 rwl_27_7 rwl_27_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_8 rbl_26_8 rbl_27_8 rc_unit R0=Rrbl C0=Crbl
xgc_27_9 wwl_27_9 wbl_27_9 rwl_27_9 rbl_27_9 sn_27_9 wos_ros_gc
xrc_wwl_27_9 wwl_27_8 wwl_27_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_9 wbl_26_9 wbl_27_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_9 rwl_27_8 rwl_27_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_9 rbl_26_9 rbl_27_9 rc_unit R0=Rrbl C0=Crbl
xgc_27_10 wwl_27_10 wbl_27_10 rwl_27_10 rbl_27_10 sn_27_10 wos_ros_gc
xrc_wwl_27_10 wwl_27_9 wwl_27_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_10 wbl_26_10 wbl_27_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_10 rwl_27_9 rwl_27_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_10 rbl_26_10 rbl_27_10 rc_unit R0=Rrbl C0=Crbl
xgc_27_11 wwl_27_11 wbl_27_11 rwl_27_11 rbl_27_11 sn_27_11 wos_ros_gc
xrc_wwl_27_11 wwl_27_10 wwl_27_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_11 wbl_26_11 wbl_27_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_11 rwl_27_10 rwl_27_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_11 rbl_26_11 rbl_27_11 rc_unit R0=Rrbl C0=Crbl
xgc_27_12 wwl_27_12 wbl_27_12 rwl_27_12 rbl_27_12 sn_27_12 wos_ros_gc
xrc_wwl_27_12 wwl_27_11 wwl_27_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_12 wbl_26_12 wbl_27_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_12 rwl_27_11 rwl_27_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_12 rbl_26_12 rbl_27_12 rc_unit R0=Rrbl C0=Crbl
xgc_27_13 wwl_27_13 wbl_27_13 rwl_27_13 rbl_27_13 sn_27_13 wos_ros_gc
xrc_wwl_27_13 wwl_27_12 wwl_27_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_13 wbl_26_13 wbl_27_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_13 rwl_27_12 rwl_27_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_13 rbl_26_13 rbl_27_13 rc_unit R0=Rrbl C0=Crbl
xgc_27_14 wwl_27_14 wbl_27_14 rwl_27_14 rbl_27_14 sn_27_14 wos_ros_gc
xrc_wwl_27_14 wwl_27_13 wwl_27_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_14 wbl_26_14 wbl_27_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_14 rwl_27_13 rwl_27_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_14 rbl_26_14 rbl_27_14 rc_unit R0=Rrbl C0=Crbl
xgc_27_15 wwl_27_15 wbl_27_15 rwl_27_15 rbl_27_15 sn_27_15 wos_ros_gc
xrc_wwl_27_15 wwl_27_14 wwl_27_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_15 wbl_26_15 wbl_27_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_15 rwl_27_14 rwl_27_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_15 rbl_26_15 rbl_27_15 rc_unit R0=Rrbl C0=Crbl
xgc_27_16 wwl_27_16 wbl_27_16 rwl_27_16 rbl_27_16 sn_27_16 wos_ros_gc
xrc_wwl_27_16 wwl_27_15 wwl_27_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_16 wbl_26_16 wbl_27_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_16 rwl_27_15 rwl_27_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_16 rbl_26_16 rbl_27_16 rc_unit R0=Rrbl C0=Crbl
xgc_27_17 wwl_27_17 wbl_27_17 rwl_27_17 rbl_27_17 sn_27_17 wos_ros_gc
xrc_wwl_27_17 wwl_27_16 wwl_27_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_17 wbl_26_17 wbl_27_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_17 rwl_27_16 rwl_27_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_17 rbl_26_17 rbl_27_17 rc_unit R0=Rrbl C0=Crbl
xgc_27_18 wwl_27_18 wbl_27_18 rwl_27_18 rbl_27_18 sn_27_18 wos_ros_gc
xrc_wwl_27_18 wwl_27_17 wwl_27_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_18 wbl_26_18 wbl_27_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_18 rwl_27_17 rwl_27_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_18 rbl_26_18 rbl_27_18 rc_unit R0=Rrbl C0=Crbl
xgc_27_19 wwl_27_19 wbl_27_19 rwl_27_19 rbl_27_19 sn_27_19 wos_ros_gc
xrc_wwl_27_19 wwl_27_18 wwl_27_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_19 wbl_26_19 wbl_27_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_19 rwl_27_18 rwl_27_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_19 rbl_26_19 rbl_27_19 rc_unit R0=Rrbl C0=Crbl
xgc_27_20 wwl_27_20 wbl_27_20 rwl_27_20 rbl_27_20 sn_27_20 wos_ros_gc
xrc_wwl_27_20 wwl_27_19 wwl_27_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_20 wbl_26_20 wbl_27_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_20 rwl_27_19 rwl_27_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_20 rbl_26_20 rbl_27_20 rc_unit R0=Rrbl C0=Crbl
xgc_27_21 wwl_27_21 wbl_27_21 rwl_27_21 rbl_27_21 sn_27_21 wos_ros_gc
xrc_wwl_27_21 wwl_27_20 wwl_27_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_21 wbl_26_21 wbl_27_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_21 rwl_27_20 rwl_27_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_21 rbl_26_21 rbl_27_21 rc_unit R0=Rrbl C0=Crbl
xgc_27_22 wwl_27_22 wbl_27_22 rwl_27_22 rbl_27_22 sn_27_22 wos_ros_gc
xrc_wwl_27_22 wwl_27_21 wwl_27_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_22 wbl_26_22 wbl_27_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_22 rwl_27_21 rwl_27_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_22 rbl_26_22 rbl_27_22 rc_unit R0=Rrbl C0=Crbl
xgc_27_23 wwl_27_23 wbl_27_23 rwl_27_23 rbl_27_23 sn_27_23 wos_ros_gc
xrc_wwl_27_23 wwl_27_22 wwl_27_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_23 wbl_26_23 wbl_27_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_23 rwl_27_22 rwl_27_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_23 rbl_26_23 rbl_27_23 rc_unit R0=Rrbl C0=Crbl
xgc_27_24 wwl_27_24 wbl_27_24 rwl_27_24 rbl_27_24 sn_27_24 wos_ros_gc
xrc_wwl_27_24 wwl_27_23 wwl_27_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_24 wbl_26_24 wbl_27_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_24 rwl_27_23 rwl_27_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_24 rbl_26_24 rbl_27_24 rc_unit R0=Rrbl C0=Crbl
xgc_27_25 wwl_27_25 wbl_27_25 rwl_27_25 rbl_27_25 sn_27_25 wos_ros_gc
xrc_wwl_27_25 wwl_27_24 wwl_27_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_25 wbl_26_25 wbl_27_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_25 rwl_27_24 rwl_27_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_25 rbl_26_25 rbl_27_25 rc_unit R0=Rrbl C0=Crbl
xgc_27_26 wwl_27_26 wbl_27_26 rwl_27_26 rbl_27_26 sn_27_26 wos_ros_gc
xrc_wwl_27_26 wwl_27_25 wwl_27_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_26 wbl_26_26 wbl_27_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_26 rwl_27_25 rwl_27_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_26 rbl_26_26 rbl_27_26 rc_unit R0=Rrbl C0=Crbl
xgc_27_27 wwl_27_27 wbl_27_27 rwl_27_27 rbl_27_27 sn_27_27 wos_ros_gc
xrc_wwl_27_27 wwl_27_26 wwl_27_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_27 wbl_26_27 wbl_27_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_27 rwl_27_26 rwl_27_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_27 rbl_26_27 rbl_27_27 rc_unit R0=Rrbl C0=Crbl
xgc_27_28 wwl_27_28 wbl_27_28 rwl_27_28 rbl_27_28 sn_27_28 wos_ros_gc
xrc_wwl_27_28 wwl_27_27 wwl_27_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_28 wbl_26_28 wbl_27_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_28 rwl_27_27 rwl_27_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_28 rbl_26_28 rbl_27_28 rc_unit R0=Rrbl C0=Crbl
xgc_27_29 wwl_27_29 wbl_27_29 rwl_27_29 rbl_27_29 sn_27_29 wos_ros_gc
xrc_wwl_27_29 wwl_27_28 wwl_27_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_29 wbl_26_29 wbl_27_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_29 rwl_27_28 rwl_27_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_29 rbl_26_29 rbl_27_29 rc_unit R0=Rrbl C0=Crbl
xgc_27_30 wwl_27_30 wbl_27_30 rwl_27_30 rbl_27_30 sn_27_30 wos_ros_gc
xrc_wwl_27_30 wwl_27_29 wwl_27_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_30 wbl_26_30 wbl_27_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_30 rwl_27_29 rwl_27_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_30 rbl_26_30 rbl_27_30 rc_unit R0=Rrbl C0=Crbl
xgc_27_31 wwl_27_31 wbl_27_31 rwl_27_31 rbl_27_31 sn_27_31 wos_ros_gc
xrc_wwl_27_31 wwl_27_30 wwl_27_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_27_31 wbl_26_31 wbl_27_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_27_31 rwl_27_30 rwl_27_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_27_31 rbl_26_31 rbl_27_31 rc_unit R0=Rrbl C0=Crbl
xgc_28_0 wwl_28_0 wbl_28_0 rwl_28_0 rbl_28_0 sn_28_0 wos_ros_gc
xrc_wwl_28_0 wwl_28 wwl_28_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_0 wbl_27_0 wbl_28_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_0 rwl_28 rwl_28_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_0 rbl_27_0 rbl_28_0 rc_unit R0=Rrbl C0=Crbl
xgc_28_1 wwl_28_1 wbl_28_1 rwl_28_1 rbl_28_1 sn_28_1 wos_ros_gc
xrc_wwl_28_1 wwl_28_0 wwl_28_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_1 wbl_27_1 wbl_28_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_1 rwl_28_0 rwl_28_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_1 rbl_27_1 rbl_28_1 rc_unit R0=Rrbl C0=Crbl
xgc_28_2 wwl_28_2 wbl_28_2 rwl_28_2 rbl_28_2 sn_28_2 wos_ros_gc
xrc_wwl_28_2 wwl_28_1 wwl_28_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_2 wbl_27_2 wbl_28_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_2 rwl_28_1 rwl_28_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_2 rbl_27_2 rbl_28_2 rc_unit R0=Rrbl C0=Crbl
xgc_28_3 wwl_28_3 wbl_28_3 rwl_28_3 rbl_28_3 sn_28_3 wos_ros_gc
xrc_wwl_28_3 wwl_28_2 wwl_28_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_3 wbl_27_3 wbl_28_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_3 rwl_28_2 rwl_28_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_3 rbl_27_3 rbl_28_3 rc_unit R0=Rrbl C0=Crbl
xgc_28_4 wwl_28_4 wbl_28_4 rwl_28_4 rbl_28_4 sn_28_4 wos_ros_gc
xrc_wwl_28_4 wwl_28_3 wwl_28_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_4 wbl_27_4 wbl_28_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_4 rwl_28_3 rwl_28_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_4 rbl_27_4 rbl_28_4 rc_unit R0=Rrbl C0=Crbl
xgc_28_5 wwl_28_5 wbl_28_5 rwl_28_5 rbl_28_5 sn_28_5 wos_ros_gc
xrc_wwl_28_5 wwl_28_4 wwl_28_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_5 wbl_27_5 wbl_28_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_5 rwl_28_4 rwl_28_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_5 rbl_27_5 rbl_28_5 rc_unit R0=Rrbl C0=Crbl
xgc_28_6 wwl_28_6 wbl_28_6 rwl_28_6 rbl_28_6 sn_28_6 wos_ros_gc
xrc_wwl_28_6 wwl_28_5 wwl_28_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_6 wbl_27_6 wbl_28_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_6 rwl_28_5 rwl_28_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_6 rbl_27_6 rbl_28_6 rc_unit R0=Rrbl C0=Crbl
xgc_28_7 wwl_28_7 wbl_28_7 rwl_28_7 rbl_28_7 sn_28_7 wos_ros_gc
xrc_wwl_28_7 wwl_28_6 wwl_28_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_7 wbl_27_7 wbl_28_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_7 rwl_28_6 rwl_28_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_7 rbl_27_7 rbl_28_7 rc_unit R0=Rrbl C0=Crbl
xgc_28_8 wwl_28_8 wbl_28_8 rwl_28_8 rbl_28_8 sn_28_8 wos_ros_gc
xrc_wwl_28_8 wwl_28_7 wwl_28_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_8 wbl_27_8 wbl_28_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_8 rwl_28_7 rwl_28_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_8 rbl_27_8 rbl_28_8 rc_unit R0=Rrbl C0=Crbl
xgc_28_9 wwl_28_9 wbl_28_9 rwl_28_9 rbl_28_9 sn_28_9 wos_ros_gc
xrc_wwl_28_9 wwl_28_8 wwl_28_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_9 wbl_27_9 wbl_28_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_9 rwl_28_8 rwl_28_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_9 rbl_27_9 rbl_28_9 rc_unit R0=Rrbl C0=Crbl
xgc_28_10 wwl_28_10 wbl_28_10 rwl_28_10 rbl_28_10 sn_28_10 wos_ros_gc
xrc_wwl_28_10 wwl_28_9 wwl_28_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_10 wbl_27_10 wbl_28_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_10 rwl_28_9 rwl_28_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_10 rbl_27_10 rbl_28_10 rc_unit R0=Rrbl C0=Crbl
xgc_28_11 wwl_28_11 wbl_28_11 rwl_28_11 rbl_28_11 sn_28_11 wos_ros_gc
xrc_wwl_28_11 wwl_28_10 wwl_28_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_11 wbl_27_11 wbl_28_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_11 rwl_28_10 rwl_28_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_11 rbl_27_11 rbl_28_11 rc_unit R0=Rrbl C0=Crbl
xgc_28_12 wwl_28_12 wbl_28_12 rwl_28_12 rbl_28_12 sn_28_12 wos_ros_gc
xrc_wwl_28_12 wwl_28_11 wwl_28_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_12 wbl_27_12 wbl_28_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_12 rwl_28_11 rwl_28_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_12 rbl_27_12 rbl_28_12 rc_unit R0=Rrbl C0=Crbl
xgc_28_13 wwl_28_13 wbl_28_13 rwl_28_13 rbl_28_13 sn_28_13 wos_ros_gc
xrc_wwl_28_13 wwl_28_12 wwl_28_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_13 wbl_27_13 wbl_28_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_13 rwl_28_12 rwl_28_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_13 rbl_27_13 rbl_28_13 rc_unit R0=Rrbl C0=Crbl
xgc_28_14 wwl_28_14 wbl_28_14 rwl_28_14 rbl_28_14 sn_28_14 wos_ros_gc
xrc_wwl_28_14 wwl_28_13 wwl_28_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_14 wbl_27_14 wbl_28_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_14 rwl_28_13 rwl_28_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_14 rbl_27_14 rbl_28_14 rc_unit R0=Rrbl C0=Crbl
xgc_28_15 wwl_28_15 wbl_28_15 rwl_28_15 rbl_28_15 sn_28_15 wos_ros_gc
xrc_wwl_28_15 wwl_28_14 wwl_28_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_15 wbl_27_15 wbl_28_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_15 rwl_28_14 rwl_28_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_15 rbl_27_15 rbl_28_15 rc_unit R0=Rrbl C0=Crbl
xgc_28_16 wwl_28_16 wbl_28_16 rwl_28_16 rbl_28_16 sn_28_16 wos_ros_gc
xrc_wwl_28_16 wwl_28_15 wwl_28_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_16 wbl_27_16 wbl_28_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_16 rwl_28_15 rwl_28_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_16 rbl_27_16 rbl_28_16 rc_unit R0=Rrbl C0=Crbl
xgc_28_17 wwl_28_17 wbl_28_17 rwl_28_17 rbl_28_17 sn_28_17 wos_ros_gc
xrc_wwl_28_17 wwl_28_16 wwl_28_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_17 wbl_27_17 wbl_28_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_17 rwl_28_16 rwl_28_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_17 rbl_27_17 rbl_28_17 rc_unit R0=Rrbl C0=Crbl
xgc_28_18 wwl_28_18 wbl_28_18 rwl_28_18 rbl_28_18 sn_28_18 wos_ros_gc
xrc_wwl_28_18 wwl_28_17 wwl_28_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_18 wbl_27_18 wbl_28_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_18 rwl_28_17 rwl_28_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_18 rbl_27_18 rbl_28_18 rc_unit R0=Rrbl C0=Crbl
xgc_28_19 wwl_28_19 wbl_28_19 rwl_28_19 rbl_28_19 sn_28_19 wos_ros_gc
xrc_wwl_28_19 wwl_28_18 wwl_28_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_19 wbl_27_19 wbl_28_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_19 rwl_28_18 rwl_28_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_19 rbl_27_19 rbl_28_19 rc_unit R0=Rrbl C0=Crbl
xgc_28_20 wwl_28_20 wbl_28_20 rwl_28_20 rbl_28_20 sn_28_20 wos_ros_gc
xrc_wwl_28_20 wwl_28_19 wwl_28_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_20 wbl_27_20 wbl_28_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_20 rwl_28_19 rwl_28_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_20 rbl_27_20 rbl_28_20 rc_unit R0=Rrbl C0=Crbl
xgc_28_21 wwl_28_21 wbl_28_21 rwl_28_21 rbl_28_21 sn_28_21 wos_ros_gc
xrc_wwl_28_21 wwl_28_20 wwl_28_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_21 wbl_27_21 wbl_28_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_21 rwl_28_20 rwl_28_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_21 rbl_27_21 rbl_28_21 rc_unit R0=Rrbl C0=Crbl
xgc_28_22 wwl_28_22 wbl_28_22 rwl_28_22 rbl_28_22 sn_28_22 wos_ros_gc
xrc_wwl_28_22 wwl_28_21 wwl_28_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_22 wbl_27_22 wbl_28_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_22 rwl_28_21 rwl_28_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_22 rbl_27_22 rbl_28_22 rc_unit R0=Rrbl C0=Crbl
xgc_28_23 wwl_28_23 wbl_28_23 rwl_28_23 rbl_28_23 sn_28_23 wos_ros_gc
xrc_wwl_28_23 wwl_28_22 wwl_28_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_23 wbl_27_23 wbl_28_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_23 rwl_28_22 rwl_28_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_23 rbl_27_23 rbl_28_23 rc_unit R0=Rrbl C0=Crbl
xgc_28_24 wwl_28_24 wbl_28_24 rwl_28_24 rbl_28_24 sn_28_24 wos_ros_gc
xrc_wwl_28_24 wwl_28_23 wwl_28_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_24 wbl_27_24 wbl_28_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_24 rwl_28_23 rwl_28_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_24 rbl_27_24 rbl_28_24 rc_unit R0=Rrbl C0=Crbl
xgc_28_25 wwl_28_25 wbl_28_25 rwl_28_25 rbl_28_25 sn_28_25 wos_ros_gc
xrc_wwl_28_25 wwl_28_24 wwl_28_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_25 wbl_27_25 wbl_28_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_25 rwl_28_24 rwl_28_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_25 rbl_27_25 rbl_28_25 rc_unit R0=Rrbl C0=Crbl
xgc_28_26 wwl_28_26 wbl_28_26 rwl_28_26 rbl_28_26 sn_28_26 wos_ros_gc
xrc_wwl_28_26 wwl_28_25 wwl_28_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_26 wbl_27_26 wbl_28_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_26 rwl_28_25 rwl_28_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_26 rbl_27_26 rbl_28_26 rc_unit R0=Rrbl C0=Crbl
xgc_28_27 wwl_28_27 wbl_28_27 rwl_28_27 rbl_28_27 sn_28_27 wos_ros_gc
xrc_wwl_28_27 wwl_28_26 wwl_28_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_27 wbl_27_27 wbl_28_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_27 rwl_28_26 rwl_28_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_27 rbl_27_27 rbl_28_27 rc_unit R0=Rrbl C0=Crbl
xgc_28_28 wwl_28_28 wbl_28_28 rwl_28_28 rbl_28_28 sn_28_28 wos_ros_gc
xrc_wwl_28_28 wwl_28_27 wwl_28_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_28 wbl_27_28 wbl_28_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_28 rwl_28_27 rwl_28_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_28 rbl_27_28 rbl_28_28 rc_unit R0=Rrbl C0=Crbl
xgc_28_29 wwl_28_29 wbl_28_29 rwl_28_29 rbl_28_29 sn_28_29 wos_ros_gc
xrc_wwl_28_29 wwl_28_28 wwl_28_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_29 wbl_27_29 wbl_28_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_29 rwl_28_28 rwl_28_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_29 rbl_27_29 rbl_28_29 rc_unit R0=Rrbl C0=Crbl
xgc_28_30 wwl_28_30 wbl_28_30 rwl_28_30 rbl_28_30 sn_28_30 wos_ros_gc
xrc_wwl_28_30 wwl_28_29 wwl_28_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_30 wbl_27_30 wbl_28_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_30 rwl_28_29 rwl_28_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_30 rbl_27_30 rbl_28_30 rc_unit R0=Rrbl C0=Crbl
xgc_28_31 wwl_28_31 wbl_28_31 rwl_28_31 rbl_28_31 sn_28_31 wos_ros_gc
xrc_wwl_28_31 wwl_28_30 wwl_28_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_28_31 wbl_27_31 wbl_28_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_28_31 rwl_28_30 rwl_28_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_28_31 rbl_27_31 rbl_28_31 rc_unit R0=Rrbl C0=Crbl
xgc_29_0 wwl_29_0 wbl_29_0 rwl_29_0 rbl_29_0 sn_29_0 wos_ros_gc
xrc_wwl_29_0 wwl_29 wwl_29_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_0 wbl_28_0 wbl_29_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_0 rwl_29 rwl_29_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_0 rbl_28_0 rbl_29_0 rc_unit R0=Rrbl C0=Crbl
xgc_29_1 wwl_29_1 wbl_29_1 rwl_29_1 rbl_29_1 sn_29_1 wos_ros_gc
xrc_wwl_29_1 wwl_29_0 wwl_29_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_1 wbl_28_1 wbl_29_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_1 rwl_29_0 rwl_29_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_1 rbl_28_1 rbl_29_1 rc_unit R0=Rrbl C0=Crbl
xgc_29_2 wwl_29_2 wbl_29_2 rwl_29_2 rbl_29_2 sn_29_2 wos_ros_gc
xrc_wwl_29_2 wwl_29_1 wwl_29_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_2 wbl_28_2 wbl_29_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_2 rwl_29_1 rwl_29_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_2 rbl_28_2 rbl_29_2 rc_unit R0=Rrbl C0=Crbl
xgc_29_3 wwl_29_3 wbl_29_3 rwl_29_3 rbl_29_3 sn_29_3 wos_ros_gc
xrc_wwl_29_3 wwl_29_2 wwl_29_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_3 wbl_28_3 wbl_29_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_3 rwl_29_2 rwl_29_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_3 rbl_28_3 rbl_29_3 rc_unit R0=Rrbl C0=Crbl
xgc_29_4 wwl_29_4 wbl_29_4 rwl_29_4 rbl_29_4 sn_29_4 wos_ros_gc
xrc_wwl_29_4 wwl_29_3 wwl_29_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_4 wbl_28_4 wbl_29_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_4 rwl_29_3 rwl_29_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_4 rbl_28_4 rbl_29_4 rc_unit R0=Rrbl C0=Crbl
xgc_29_5 wwl_29_5 wbl_29_5 rwl_29_5 rbl_29_5 sn_29_5 wos_ros_gc
xrc_wwl_29_5 wwl_29_4 wwl_29_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_5 wbl_28_5 wbl_29_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_5 rwl_29_4 rwl_29_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_5 rbl_28_5 rbl_29_5 rc_unit R0=Rrbl C0=Crbl
xgc_29_6 wwl_29_6 wbl_29_6 rwl_29_6 rbl_29_6 sn_29_6 wos_ros_gc
xrc_wwl_29_6 wwl_29_5 wwl_29_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_6 wbl_28_6 wbl_29_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_6 rwl_29_5 rwl_29_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_6 rbl_28_6 rbl_29_6 rc_unit R0=Rrbl C0=Crbl
xgc_29_7 wwl_29_7 wbl_29_7 rwl_29_7 rbl_29_7 sn_29_7 wos_ros_gc
xrc_wwl_29_7 wwl_29_6 wwl_29_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_7 wbl_28_7 wbl_29_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_7 rwl_29_6 rwl_29_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_7 rbl_28_7 rbl_29_7 rc_unit R0=Rrbl C0=Crbl
xgc_29_8 wwl_29_8 wbl_29_8 rwl_29_8 rbl_29_8 sn_29_8 wos_ros_gc
xrc_wwl_29_8 wwl_29_7 wwl_29_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_8 wbl_28_8 wbl_29_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_8 rwl_29_7 rwl_29_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_8 rbl_28_8 rbl_29_8 rc_unit R0=Rrbl C0=Crbl
xgc_29_9 wwl_29_9 wbl_29_9 rwl_29_9 rbl_29_9 sn_29_9 wos_ros_gc
xrc_wwl_29_9 wwl_29_8 wwl_29_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_9 wbl_28_9 wbl_29_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_9 rwl_29_8 rwl_29_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_9 rbl_28_9 rbl_29_9 rc_unit R0=Rrbl C0=Crbl
xgc_29_10 wwl_29_10 wbl_29_10 rwl_29_10 rbl_29_10 sn_29_10 wos_ros_gc
xrc_wwl_29_10 wwl_29_9 wwl_29_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_10 wbl_28_10 wbl_29_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_10 rwl_29_9 rwl_29_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_10 rbl_28_10 rbl_29_10 rc_unit R0=Rrbl C0=Crbl
xgc_29_11 wwl_29_11 wbl_29_11 rwl_29_11 rbl_29_11 sn_29_11 wos_ros_gc
xrc_wwl_29_11 wwl_29_10 wwl_29_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_11 wbl_28_11 wbl_29_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_11 rwl_29_10 rwl_29_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_11 rbl_28_11 rbl_29_11 rc_unit R0=Rrbl C0=Crbl
xgc_29_12 wwl_29_12 wbl_29_12 rwl_29_12 rbl_29_12 sn_29_12 wos_ros_gc
xrc_wwl_29_12 wwl_29_11 wwl_29_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_12 wbl_28_12 wbl_29_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_12 rwl_29_11 rwl_29_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_12 rbl_28_12 rbl_29_12 rc_unit R0=Rrbl C0=Crbl
xgc_29_13 wwl_29_13 wbl_29_13 rwl_29_13 rbl_29_13 sn_29_13 wos_ros_gc
xrc_wwl_29_13 wwl_29_12 wwl_29_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_13 wbl_28_13 wbl_29_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_13 rwl_29_12 rwl_29_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_13 rbl_28_13 rbl_29_13 rc_unit R0=Rrbl C0=Crbl
xgc_29_14 wwl_29_14 wbl_29_14 rwl_29_14 rbl_29_14 sn_29_14 wos_ros_gc
xrc_wwl_29_14 wwl_29_13 wwl_29_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_14 wbl_28_14 wbl_29_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_14 rwl_29_13 rwl_29_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_14 rbl_28_14 rbl_29_14 rc_unit R0=Rrbl C0=Crbl
xgc_29_15 wwl_29_15 wbl_29_15 rwl_29_15 rbl_29_15 sn_29_15 wos_ros_gc
xrc_wwl_29_15 wwl_29_14 wwl_29_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_15 wbl_28_15 wbl_29_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_15 rwl_29_14 rwl_29_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_15 rbl_28_15 rbl_29_15 rc_unit R0=Rrbl C0=Crbl
xgc_29_16 wwl_29_16 wbl_29_16 rwl_29_16 rbl_29_16 sn_29_16 wos_ros_gc
xrc_wwl_29_16 wwl_29_15 wwl_29_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_16 wbl_28_16 wbl_29_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_16 rwl_29_15 rwl_29_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_16 rbl_28_16 rbl_29_16 rc_unit R0=Rrbl C0=Crbl
xgc_29_17 wwl_29_17 wbl_29_17 rwl_29_17 rbl_29_17 sn_29_17 wos_ros_gc
xrc_wwl_29_17 wwl_29_16 wwl_29_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_17 wbl_28_17 wbl_29_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_17 rwl_29_16 rwl_29_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_17 rbl_28_17 rbl_29_17 rc_unit R0=Rrbl C0=Crbl
xgc_29_18 wwl_29_18 wbl_29_18 rwl_29_18 rbl_29_18 sn_29_18 wos_ros_gc
xrc_wwl_29_18 wwl_29_17 wwl_29_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_18 wbl_28_18 wbl_29_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_18 rwl_29_17 rwl_29_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_18 rbl_28_18 rbl_29_18 rc_unit R0=Rrbl C0=Crbl
xgc_29_19 wwl_29_19 wbl_29_19 rwl_29_19 rbl_29_19 sn_29_19 wos_ros_gc
xrc_wwl_29_19 wwl_29_18 wwl_29_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_19 wbl_28_19 wbl_29_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_19 rwl_29_18 rwl_29_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_19 rbl_28_19 rbl_29_19 rc_unit R0=Rrbl C0=Crbl
xgc_29_20 wwl_29_20 wbl_29_20 rwl_29_20 rbl_29_20 sn_29_20 wos_ros_gc
xrc_wwl_29_20 wwl_29_19 wwl_29_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_20 wbl_28_20 wbl_29_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_20 rwl_29_19 rwl_29_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_20 rbl_28_20 rbl_29_20 rc_unit R0=Rrbl C0=Crbl
xgc_29_21 wwl_29_21 wbl_29_21 rwl_29_21 rbl_29_21 sn_29_21 wos_ros_gc
xrc_wwl_29_21 wwl_29_20 wwl_29_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_21 wbl_28_21 wbl_29_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_21 rwl_29_20 rwl_29_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_21 rbl_28_21 rbl_29_21 rc_unit R0=Rrbl C0=Crbl
xgc_29_22 wwl_29_22 wbl_29_22 rwl_29_22 rbl_29_22 sn_29_22 wos_ros_gc
xrc_wwl_29_22 wwl_29_21 wwl_29_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_22 wbl_28_22 wbl_29_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_22 rwl_29_21 rwl_29_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_22 rbl_28_22 rbl_29_22 rc_unit R0=Rrbl C0=Crbl
xgc_29_23 wwl_29_23 wbl_29_23 rwl_29_23 rbl_29_23 sn_29_23 wos_ros_gc
xrc_wwl_29_23 wwl_29_22 wwl_29_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_23 wbl_28_23 wbl_29_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_23 rwl_29_22 rwl_29_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_23 rbl_28_23 rbl_29_23 rc_unit R0=Rrbl C0=Crbl
xgc_29_24 wwl_29_24 wbl_29_24 rwl_29_24 rbl_29_24 sn_29_24 wos_ros_gc
xrc_wwl_29_24 wwl_29_23 wwl_29_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_24 wbl_28_24 wbl_29_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_24 rwl_29_23 rwl_29_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_24 rbl_28_24 rbl_29_24 rc_unit R0=Rrbl C0=Crbl
xgc_29_25 wwl_29_25 wbl_29_25 rwl_29_25 rbl_29_25 sn_29_25 wos_ros_gc
xrc_wwl_29_25 wwl_29_24 wwl_29_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_25 wbl_28_25 wbl_29_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_25 rwl_29_24 rwl_29_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_25 rbl_28_25 rbl_29_25 rc_unit R0=Rrbl C0=Crbl
xgc_29_26 wwl_29_26 wbl_29_26 rwl_29_26 rbl_29_26 sn_29_26 wos_ros_gc
xrc_wwl_29_26 wwl_29_25 wwl_29_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_26 wbl_28_26 wbl_29_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_26 rwl_29_25 rwl_29_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_26 rbl_28_26 rbl_29_26 rc_unit R0=Rrbl C0=Crbl
xgc_29_27 wwl_29_27 wbl_29_27 rwl_29_27 rbl_29_27 sn_29_27 wos_ros_gc
xrc_wwl_29_27 wwl_29_26 wwl_29_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_27 wbl_28_27 wbl_29_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_27 rwl_29_26 rwl_29_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_27 rbl_28_27 rbl_29_27 rc_unit R0=Rrbl C0=Crbl
xgc_29_28 wwl_29_28 wbl_29_28 rwl_29_28 rbl_29_28 sn_29_28 wos_ros_gc
xrc_wwl_29_28 wwl_29_27 wwl_29_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_28 wbl_28_28 wbl_29_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_28 rwl_29_27 rwl_29_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_28 rbl_28_28 rbl_29_28 rc_unit R0=Rrbl C0=Crbl
xgc_29_29 wwl_29_29 wbl_29_29 rwl_29_29 rbl_29_29 sn_29_29 wos_ros_gc
xrc_wwl_29_29 wwl_29_28 wwl_29_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_29 wbl_28_29 wbl_29_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_29 rwl_29_28 rwl_29_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_29 rbl_28_29 rbl_29_29 rc_unit R0=Rrbl C0=Crbl
xgc_29_30 wwl_29_30 wbl_29_30 rwl_29_30 rbl_29_30 sn_29_30 wos_ros_gc
xrc_wwl_29_30 wwl_29_29 wwl_29_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_30 wbl_28_30 wbl_29_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_30 rwl_29_29 rwl_29_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_30 rbl_28_30 rbl_29_30 rc_unit R0=Rrbl C0=Crbl
xgc_29_31 wwl_29_31 wbl_29_31 rwl_29_31 rbl_29_31 sn_29_31 wos_ros_gc
xrc_wwl_29_31 wwl_29_30 wwl_29_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_29_31 wbl_28_31 wbl_29_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_29_31 rwl_29_30 rwl_29_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_29_31 rbl_28_31 rbl_29_31 rc_unit R0=Rrbl C0=Crbl
xgc_30_0 wwl_30_0 wbl_30_0 rwl_30_0 rbl_30_0 sn_30_0 wos_ros_gc
xrc_wwl_30_0 wwl_30 wwl_30_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_0 wbl_29_0 wbl_30_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_0 rwl_30 rwl_30_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_0 rbl_29_0 rbl_30_0 rc_unit R0=Rrbl C0=Crbl
xgc_30_1 wwl_30_1 wbl_30_1 rwl_30_1 rbl_30_1 sn_30_1 wos_ros_gc
xrc_wwl_30_1 wwl_30_0 wwl_30_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_1 wbl_29_1 wbl_30_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_1 rwl_30_0 rwl_30_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_1 rbl_29_1 rbl_30_1 rc_unit R0=Rrbl C0=Crbl
xgc_30_2 wwl_30_2 wbl_30_2 rwl_30_2 rbl_30_2 sn_30_2 wos_ros_gc
xrc_wwl_30_2 wwl_30_1 wwl_30_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_2 wbl_29_2 wbl_30_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_2 rwl_30_1 rwl_30_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_2 rbl_29_2 rbl_30_2 rc_unit R0=Rrbl C0=Crbl
xgc_30_3 wwl_30_3 wbl_30_3 rwl_30_3 rbl_30_3 sn_30_3 wos_ros_gc
xrc_wwl_30_3 wwl_30_2 wwl_30_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_3 wbl_29_3 wbl_30_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_3 rwl_30_2 rwl_30_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_3 rbl_29_3 rbl_30_3 rc_unit R0=Rrbl C0=Crbl
xgc_30_4 wwl_30_4 wbl_30_4 rwl_30_4 rbl_30_4 sn_30_4 wos_ros_gc
xrc_wwl_30_4 wwl_30_3 wwl_30_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_4 wbl_29_4 wbl_30_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_4 rwl_30_3 rwl_30_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_4 rbl_29_4 rbl_30_4 rc_unit R0=Rrbl C0=Crbl
xgc_30_5 wwl_30_5 wbl_30_5 rwl_30_5 rbl_30_5 sn_30_5 wos_ros_gc
xrc_wwl_30_5 wwl_30_4 wwl_30_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_5 wbl_29_5 wbl_30_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_5 rwl_30_4 rwl_30_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_5 rbl_29_5 rbl_30_5 rc_unit R0=Rrbl C0=Crbl
xgc_30_6 wwl_30_6 wbl_30_6 rwl_30_6 rbl_30_6 sn_30_6 wos_ros_gc
xrc_wwl_30_6 wwl_30_5 wwl_30_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_6 wbl_29_6 wbl_30_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_6 rwl_30_5 rwl_30_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_6 rbl_29_6 rbl_30_6 rc_unit R0=Rrbl C0=Crbl
xgc_30_7 wwl_30_7 wbl_30_7 rwl_30_7 rbl_30_7 sn_30_7 wos_ros_gc
xrc_wwl_30_7 wwl_30_6 wwl_30_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_7 wbl_29_7 wbl_30_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_7 rwl_30_6 rwl_30_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_7 rbl_29_7 rbl_30_7 rc_unit R0=Rrbl C0=Crbl
xgc_30_8 wwl_30_8 wbl_30_8 rwl_30_8 rbl_30_8 sn_30_8 wos_ros_gc
xrc_wwl_30_8 wwl_30_7 wwl_30_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_8 wbl_29_8 wbl_30_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_8 rwl_30_7 rwl_30_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_8 rbl_29_8 rbl_30_8 rc_unit R0=Rrbl C0=Crbl
xgc_30_9 wwl_30_9 wbl_30_9 rwl_30_9 rbl_30_9 sn_30_9 wos_ros_gc
xrc_wwl_30_9 wwl_30_8 wwl_30_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_9 wbl_29_9 wbl_30_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_9 rwl_30_8 rwl_30_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_9 rbl_29_9 rbl_30_9 rc_unit R0=Rrbl C0=Crbl
xgc_30_10 wwl_30_10 wbl_30_10 rwl_30_10 rbl_30_10 sn_30_10 wos_ros_gc
xrc_wwl_30_10 wwl_30_9 wwl_30_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_10 wbl_29_10 wbl_30_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_10 rwl_30_9 rwl_30_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_10 rbl_29_10 rbl_30_10 rc_unit R0=Rrbl C0=Crbl
xgc_30_11 wwl_30_11 wbl_30_11 rwl_30_11 rbl_30_11 sn_30_11 wos_ros_gc
xrc_wwl_30_11 wwl_30_10 wwl_30_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_11 wbl_29_11 wbl_30_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_11 rwl_30_10 rwl_30_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_11 rbl_29_11 rbl_30_11 rc_unit R0=Rrbl C0=Crbl
xgc_30_12 wwl_30_12 wbl_30_12 rwl_30_12 rbl_30_12 sn_30_12 wos_ros_gc
xrc_wwl_30_12 wwl_30_11 wwl_30_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_12 wbl_29_12 wbl_30_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_12 rwl_30_11 rwl_30_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_12 rbl_29_12 rbl_30_12 rc_unit R0=Rrbl C0=Crbl
xgc_30_13 wwl_30_13 wbl_30_13 rwl_30_13 rbl_30_13 sn_30_13 wos_ros_gc
xrc_wwl_30_13 wwl_30_12 wwl_30_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_13 wbl_29_13 wbl_30_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_13 rwl_30_12 rwl_30_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_13 rbl_29_13 rbl_30_13 rc_unit R0=Rrbl C0=Crbl
xgc_30_14 wwl_30_14 wbl_30_14 rwl_30_14 rbl_30_14 sn_30_14 wos_ros_gc
xrc_wwl_30_14 wwl_30_13 wwl_30_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_14 wbl_29_14 wbl_30_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_14 rwl_30_13 rwl_30_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_14 rbl_29_14 rbl_30_14 rc_unit R0=Rrbl C0=Crbl
xgc_30_15 wwl_30_15 wbl_30_15 rwl_30_15 rbl_30_15 sn_30_15 wos_ros_gc
xrc_wwl_30_15 wwl_30_14 wwl_30_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_15 wbl_29_15 wbl_30_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_15 rwl_30_14 rwl_30_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_15 rbl_29_15 rbl_30_15 rc_unit R0=Rrbl C0=Crbl
xgc_30_16 wwl_30_16 wbl_30_16 rwl_30_16 rbl_30_16 sn_30_16 wos_ros_gc
xrc_wwl_30_16 wwl_30_15 wwl_30_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_16 wbl_29_16 wbl_30_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_16 rwl_30_15 rwl_30_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_16 rbl_29_16 rbl_30_16 rc_unit R0=Rrbl C0=Crbl
xgc_30_17 wwl_30_17 wbl_30_17 rwl_30_17 rbl_30_17 sn_30_17 wos_ros_gc
xrc_wwl_30_17 wwl_30_16 wwl_30_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_17 wbl_29_17 wbl_30_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_17 rwl_30_16 rwl_30_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_17 rbl_29_17 rbl_30_17 rc_unit R0=Rrbl C0=Crbl
xgc_30_18 wwl_30_18 wbl_30_18 rwl_30_18 rbl_30_18 sn_30_18 wos_ros_gc
xrc_wwl_30_18 wwl_30_17 wwl_30_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_18 wbl_29_18 wbl_30_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_18 rwl_30_17 rwl_30_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_18 rbl_29_18 rbl_30_18 rc_unit R0=Rrbl C0=Crbl
xgc_30_19 wwl_30_19 wbl_30_19 rwl_30_19 rbl_30_19 sn_30_19 wos_ros_gc
xrc_wwl_30_19 wwl_30_18 wwl_30_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_19 wbl_29_19 wbl_30_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_19 rwl_30_18 rwl_30_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_19 rbl_29_19 rbl_30_19 rc_unit R0=Rrbl C0=Crbl
xgc_30_20 wwl_30_20 wbl_30_20 rwl_30_20 rbl_30_20 sn_30_20 wos_ros_gc
xrc_wwl_30_20 wwl_30_19 wwl_30_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_20 wbl_29_20 wbl_30_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_20 rwl_30_19 rwl_30_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_20 rbl_29_20 rbl_30_20 rc_unit R0=Rrbl C0=Crbl
xgc_30_21 wwl_30_21 wbl_30_21 rwl_30_21 rbl_30_21 sn_30_21 wos_ros_gc
xrc_wwl_30_21 wwl_30_20 wwl_30_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_21 wbl_29_21 wbl_30_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_21 rwl_30_20 rwl_30_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_21 rbl_29_21 rbl_30_21 rc_unit R0=Rrbl C0=Crbl
xgc_30_22 wwl_30_22 wbl_30_22 rwl_30_22 rbl_30_22 sn_30_22 wos_ros_gc
xrc_wwl_30_22 wwl_30_21 wwl_30_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_22 wbl_29_22 wbl_30_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_22 rwl_30_21 rwl_30_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_22 rbl_29_22 rbl_30_22 rc_unit R0=Rrbl C0=Crbl
xgc_30_23 wwl_30_23 wbl_30_23 rwl_30_23 rbl_30_23 sn_30_23 wos_ros_gc
xrc_wwl_30_23 wwl_30_22 wwl_30_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_23 wbl_29_23 wbl_30_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_23 rwl_30_22 rwl_30_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_23 rbl_29_23 rbl_30_23 rc_unit R0=Rrbl C0=Crbl
xgc_30_24 wwl_30_24 wbl_30_24 rwl_30_24 rbl_30_24 sn_30_24 wos_ros_gc
xrc_wwl_30_24 wwl_30_23 wwl_30_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_24 wbl_29_24 wbl_30_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_24 rwl_30_23 rwl_30_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_24 rbl_29_24 rbl_30_24 rc_unit R0=Rrbl C0=Crbl
xgc_30_25 wwl_30_25 wbl_30_25 rwl_30_25 rbl_30_25 sn_30_25 wos_ros_gc
xrc_wwl_30_25 wwl_30_24 wwl_30_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_25 wbl_29_25 wbl_30_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_25 rwl_30_24 rwl_30_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_25 rbl_29_25 rbl_30_25 rc_unit R0=Rrbl C0=Crbl
xgc_30_26 wwl_30_26 wbl_30_26 rwl_30_26 rbl_30_26 sn_30_26 wos_ros_gc
xrc_wwl_30_26 wwl_30_25 wwl_30_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_26 wbl_29_26 wbl_30_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_26 rwl_30_25 rwl_30_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_26 rbl_29_26 rbl_30_26 rc_unit R0=Rrbl C0=Crbl
xgc_30_27 wwl_30_27 wbl_30_27 rwl_30_27 rbl_30_27 sn_30_27 wos_ros_gc
xrc_wwl_30_27 wwl_30_26 wwl_30_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_27 wbl_29_27 wbl_30_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_27 rwl_30_26 rwl_30_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_27 rbl_29_27 rbl_30_27 rc_unit R0=Rrbl C0=Crbl
xgc_30_28 wwl_30_28 wbl_30_28 rwl_30_28 rbl_30_28 sn_30_28 wos_ros_gc
xrc_wwl_30_28 wwl_30_27 wwl_30_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_28 wbl_29_28 wbl_30_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_28 rwl_30_27 rwl_30_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_28 rbl_29_28 rbl_30_28 rc_unit R0=Rrbl C0=Crbl
xgc_30_29 wwl_30_29 wbl_30_29 rwl_30_29 rbl_30_29 sn_30_29 wos_ros_gc
xrc_wwl_30_29 wwl_30_28 wwl_30_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_29 wbl_29_29 wbl_30_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_29 rwl_30_28 rwl_30_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_29 rbl_29_29 rbl_30_29 rc_unit R0=Rrbl C0=Crbl
xgc_30_30 wwl_30_30 wbl_30_30 rwl_30_30 rbl_30_30 sn_30_30 wos_ros_gc
xrc_wwl_30_30 wwl_30_29 wwl_30_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_30 wbl_29_30 wbl_30_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_30 rwl_30_29 rwl_30_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_30 rbl_29_30 rbl_30_30 rc_unit R0=Rrbl C0=Crbl
xgc_30_31 wwl_30_31 wbl_30_31 rwl_30_31 rbl_30_31 sn_30_31 wos_ros_gc
xrc_wwl_30_31 wwl_30_30 wwl_30_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_30_31 wbl_29_31 wbl_30_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_30_31 rwl_30_30 rwl_30_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_30_31 rbl_29_31 rbl_30_31 rc_unit R0=Rrbl C0=Crbl
xgc_31_0 wwl_31_0 wbl_31_0 rwl_31_0 rbl_31_0 sn_31_0 wos_ros_gc
xrc_wwl_31_0 wwl_31 wwl_31_0 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_0 wbl_30_0 wbl_31_0 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_0 rwl_31 rwl_31_0 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_0 rbl_30_0 rbl_31_0 rc_unit R0=Rrbl C0=Crbl
xgc_31_1 wwl_31_1 wbl_31_1 rwl_31_1 rbl_31_1 sn_31_1 wos_ros_gc
xrc_wwl_31_1 wwl_31_0 wwl_31_1 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_1 wbl_30_1 wbl_31_1 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_1 rwl_31_0 rwl_31_1 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_1 rbl_30_1 rbl_31_1 rc_unit R0=Rrbl C0=Crbl
xgc_31_2 wwl_31_2 wbl_31_2 rwl_31_2 rbl_31_2 sn_31_2 wos_ros_gc
xrc_wwl_31_2 wwl_31_1 wwl_31_2 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_2 wbl_30_2 wbl_31_2 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_2 rwl_31_1 rwl_31_2 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_2 rbl_30_2 rbl_31_2 rc_unit R0=Rrbl C0=Crbl
xgc_31_3 wwl_31_3 wbl_31_3 rwl_31_3 rbl_31_3 sn_31_3 wos_ros_gc
xrc_wwl_31_3 wwl_31_2 wwl_31_3 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_3 wbl_30_3 wbl_31_3 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_3 rwl_31_2 rwl_31_3 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_3 rbl_30_3 rbl_31_3 rc_unit R0=Rrbl C0=Crbl
xgc_31_4 wwl_31_4 wbl_31_4 rwl_31_4 rbl_31_4 sn_31_4 wos_ros_gc
xrc_wwl_31_4 wwl_31_3 wwl_31_4 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_4 wbl_30_4 wbl_31_4 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_4 rwl_31_3 rwl_31_4 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_4 rbl_30_4 rbl_31_4 rc_unit R0=Rrbl C0=Crbl
xgc_31_5 wwl_31_5 wbl_31_5 rwl_31_5 rbl_31_5 sn_31_5 wos_ros_gc
xrc_wwl_31_5 wwl_31_4 wwl_31_5 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_5 wbl_30_5 wbl_31_5 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_5 rwl_31_4 rwl_31_5 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_5 rbl_30_5 rbl_31_5 rc_unit R0=Rrbl C0=Crbl
xgc_31_6 wwl_31_6 wbl_31_6 rwl_31_6 rbl_31_6 sn_31_6 wos_ros_gc
xrc_wwl_31_6 wwl_31_5 wwl_31_6 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_6 wbl_30_6 wbl_31_6 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_6 rwl_31_5 rwl_31_6 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_6 rbl_30_6 rbl_31_6 rc_unit R0=Rrbl C0=Crbl
xgc_31_7 wwl_31_7 wbl_31_7 rwl_31_7 rbl_31_7 sn_31_7 wos_ros_gc
xrc_wwl_31_7 wwl_31_6 wwl_31_7 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_7 wbl_30_7 wbl_31_7 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_7 rwl_31_6 rwl_31_7 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_7 rbl_30_7 rbl_31_7 rc_unit R0=Rrbl C0=Crbl
xgc_31_8 wwl_31_8 wbl_31_8 rwl_31_8 rbl_31_8 sn_31_8 wos_ros_gc
xrc_wwl_31_8 wwl_31_7 wwl_31_8 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_8 wbl_30_8 wbl_31_8 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_8 rwl_31_7 rwl_31_8 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_8 rbl_30_8 rbl_31_8 rc_unit R0=Rrbl C0=Crbl
xgc_31_9 wwl_31_9 wbl_31_9 rwl_31_9 rbl_31_9 sn_31_9 wos_ros_gc
xrc_wwl_31_9 wwl_31_8 wwl_31_9 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_9 wbl_30_9 wbl_31_9 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_9 rwl_31_8 rwl_31_9 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_9 rbl_30_9 rbl_31_9 rc_unit R0=Rrbl C0=Crbl
xgc_31_10 wwl_31_10 wbl_31_10 rwl_31_10 rbl_31_10 sn_31_10 wos_ros_gc
xrc_wwl_31_10 wwl_31_9 wwl_31_10 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_10 wbl_30_10 wbl_31_10 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_10 rwl_31_9 rwl_31_10 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_10 rbl_30_10 rbl_31_10 rc_unit R0=Rrbl C0=Crbl
xgc_31_11 wwl_31_11 wbl_31_11 rwl_31_11 rbl_31_11 sn_31_11 wos_ros_gc
xrc_wwl_31_11 wwl_31_10 wwl_31_11 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_11 wbl_30_11 wbl_31_11 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_11 rwl_31_10 rwl_31_11 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_11 rbl_30_11 rbl_31_11 rc_unit R0=Rrbl C0=Crbl
xgc_31_12 wwl_31_12 wbl_31_12 rwl_31_12 rbl_31_12 sn_31_12 wos_ros_gc
xrc_wwl_31_12 wwl_31_11 wwl_31_12 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_12 wbl_30_12 wbl_31_12 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_12 rwl_31_11 rwl_31_12 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_12 rbl_30_12 rbl_31_12 rc_unit R0=Rrbl C0=Crbl
xgc_31_13 wwl_31_13 wbl_31_13 rwl_31_13 rbl_31_13 sn_31_13 wos_ros_gc
xrc_wwl_31_13 wwl_31_12 wwl_31_13 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_13 wbl_30_13 wbl_31_13 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_13 rwl_31_12 rwl_31_13 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_13 rbl_30_13 rbl_31_13 rc_unit R0=Rrbl C0=Crbl
xgc_31_14 wwl_31_14 wbl_31_14 rwl_31_14 rbl_31_14 sn_31_14 wos_ros_gc
xrc_wwl_31_14 wwl_31_13 wwl_31_14 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_14 wbl_30_14 wbl_31_14 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_14 rwl_31_13 rwl_31_14 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_14 rbl_30_14 rbl_31_14 rc_unit R0=Rrbl C0=Crbl
xgc_31_15 wwl_31_15 wbl_31_15 rwl_31_15 rbl_31_15 sn_31_15 wos_ros_gc
xrc_wwl_31_15 wwl_31_14 wwl_31_15 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_15 wbl_30_15 wbl_31_15 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_15 rwl_31_14 rwl_31_15 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_15 rbl_30_15 rbl_31_15 rc_unit R0=Rrbl C0=Crbl
xgc_31_16 wwl_31_16 wbl_31_16 rwl_31_16 rbl_31_16 sn_31_16 wos_ros_gc
xrc_wwl_31_16 wwl_31_15 wwl_31_16 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_16 wbl_30_16 wbl_31_16 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_16 rwl_31_15 rwl_31_16 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_16 rbl_30_16 rbl_31_16 rc_unit R0=Rrbl C0=Crbl
xgc_31_17 wwl_31_17 wbl_31_17 rwl_31_17 rbl_31_17 sn_31_17 wos_ros_gc
xrc_wwl_31_17 wwl_31_16 wwl_31_17 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_17 wbl_30_17 wbl_31_17 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_17 rwl_31_16 rwl_31_17 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_17 rbl_30_17 rbl_31_17 rc_unit R0=Rrbl C0=Crbl
xgc_31_18 wwl_31_18 wbl_31_18 rwl_31_18 rbl_31_18 sn_31_18 wos_ros_gc
xrc_wwl_31_18 wwl_31_17 wwl_31_18 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_18 wbl_30_18 wbl_31_18 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_18 rwl_31_17 rwl_31_18 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_18 rbl_30_18 rbl_31_18 rc_unit R0=Rrbl C0=Crbl
xgc_31_19 wwl_31_19 wbl_31_19 rwl_31_19 rbl_31_19 sn_31_19 wos_ros_gc
xrc_wwl_31_19 wwl_31_18 wwl_31_19 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_19 wbl_30_19 wbl_31_19 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_19 rwl_31_18 rwl_31_19 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_19 rbl_30_19 rbl_31_19 rc_unit R0=Rrbl C0=Crbl
xgc_31_20 wwl_31_20 wbl_31_20 rwl_31_20 rbl_31_20 sn_31_20 wos_ros_gc
xrc_wwl_31_20 wwl_31_19 wwl_31_20 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_20 wbl_30_20 wbl_31_20 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_20 rwl_31_19 rwl_31_20 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_20 rbl_30_20 rbl_31_20 rc_unit R0=Rrbl C0=Crbl
xgc_31_21 wwl_31_21 wbl_31_21 rwl_31_21 rbl_31_21 sn_31_21 wos_ros_gc
xrc_wwl_31_21 wwl_31_20 wwl_31_21 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_21 wbl_30_21 wbl_31_21 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_21 rwl_31_20 rwl_31_21 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_21 rbl_30_21 rbl_31_21 rc_unit R0=Rrbl C0=Crbl
xgc_31_22 wwl_31_22 wbl_31_22 rwl_31_22 rbl_31_22 sn_31_22 wos_ros_gc
xrc_wwl_31_22 wwl_31_21 wwl_31_22 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_22 wbl_30_22 wbl_31_22 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_22 rwl_31_21 rwl_31_22 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_22 rbl_30_22 rbl_31_22 rc_unit R0=Rrbl C0=Crbl
xgc_31_23 wwl_31_23 wbl_31_23 rwl_31_23 rbl_31_23 sn_31_23 wos_ros_gc
xrc_wwl_31_23 wwl_31_22 wwl_31_23 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_23 wbl_30_23 wbl_31_23 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_23 rwl_31_22 rwl_31_23 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_23 rbl_30_23 rbl_31_23 rc_unit R0=Rrbl C0=Crbl
xgc_31_24 wwl_31_24 wbl_31_24 rwl_31_24 rbl_31_24 sn_31_24 wos_ros_gc
xrc_wwl_31_24 wwl_31_23 wwl_31_24 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_24 wbl_30_24 wbl_31_24 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_24 rwl_31_23 rwl_31_24 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_24 rbl_30_24 rbl_31_24 rc_unit R0=Rrbl C0=Crbl
xgc_31_25 wwl_31_25 wbl_31_25 rwl_31_25 rbl_31_25 sn_31_25 wos_ros_gc
xrc_wwl_31_25 wwl_31_24 wwl_31_25 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_25 wbl_30_25 wbl_31_25 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_25 rwl_31_24 rwl_31_25 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_25 rbl_30_25 rbl_31_25 rc_unit R0=Rrbl C0=Crbl
xgc_31_26 wwl_31_26 wbl_31_26 rwl_31_26 rbl_31_26 sn_31_26 wos_ros_gc
xrc_wwl_31_26 wwl_31_25 wwl_31_26 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_26 wbl_30_26 wbl_31_26 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_26 rwl_31_25 rwl_31_26 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_26 rbl_30_26 rbl_31_26 rc_unit R0=Rrbl C0=Crbl
xgc_31_27 wwl_31_27 wbl_31_27 rwl_31_27 rbl_31_27 sn_31_27 wos_ros_gc
xrc_wwl_31_27 wwl_31_26 wwl_31_27 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_27 wbl_30_27 wbl_31_27 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_27 rwl_31_26 rwl_31_27 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_27 rbl_30_27 rbl_31_27 rc_unit R0=Rrbl C0=Crbl
xgc_31_28 wwl_31_28 wbl_31_28 rwl_31_28 rbl_31_28 sn_31_28 wos_ros_gc
xrc_wwl_31_28 wwl_31_27 wwl_31_28 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_28 wbl_30_28 wbl_31_28 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_28 rwl_31_27 rwl_31_28 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_28 rbl_30_28 rbl_31_28 rc_unit R0=Rrbl C0=Crbl
xgc_31_29 wwl_31_29 wbl_31_29 rwl_31_29 rbl_31_29 sn_31_29 wos_ros_gc
xrc_wwl_31_29 wwl_31_28 wwl_31_29 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_29 wbl_30_29 wbl_31_29 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_29 rwl_31_28 rwl_31_29 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_29 rbl_30_29 rbl_31_29 rc_unit R0=Rrbl C0=Crbl
xgc_31_30 wwl_31_30 wbl_31_30 rwl_31_30 rbl_31_30 sn_31_30 wos_ros_gc
xrc_wwl_31_30 wwl_31_29 wwl_31_30 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_30 wbl_30_30 wbl_31_30 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_30 rwl_31_29 rwl_31_30 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_30 rbl_30_30 rbl_31_30 rc_unit R0=Rrbl C0=Crbl
xgc_31_31 wwl_31_31 wbl_31_31 rwl_31_31 rbl_31_31 sn_31_31 wos_ros_gc
xrc_wwl_31_31 wwl_31_30 wwl_31_31 rc_unit R0=Rwwl C0=Cwwl
xrc_wbl_31_31 wbl_30_31 wbl_31_31 rc_unit R0=Rwbl C0=Cwbl
xrc_rwl_31_31 rwl_31_30 rwl_31_31 rc_unit R0=Rrwl C0=Crwl
xrc_rbl_31_31 rbl_30_31 rbl_31_31 rc_unit R0=Rrbl C0=Crbl
vww_0 wwl_0 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_0 rwl_0 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_1 wwl_1 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_1 rwl_1 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_2 wwl_2 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_2 rwl_2 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_3 wwl_3 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_3 rwl_3 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_4 wwl_4 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_4 rwl_4 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_5 wwl_5 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_5 rwl_5 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_6 wwl_6 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_6 rwl_6 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_7 wwl_7 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_7 rwl_7 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_8 wwl_8 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_8 rwl_8 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_9 wwl_9 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_9 rwl_9 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_10 wwl_10 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_10 rwl_10 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_11 wwl_11 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_11 rwl_11 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_12 wwl_12 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_12 rwl_12 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_13 wwl_13 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_13 rwl_13 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_14 wwl_14 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_14 rwl_14 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_15 wwl_15 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_15 rwl_15 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_16 wwl_16 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_16 rwl_16 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_17 wwl_17 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_17 rwl_17 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_18 wwl_18 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_18 rwl_18 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_19 wwl_19 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_19 rwl_19 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_20 wwl_20 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_20 rwl_20 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_21 wwl_21 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_21 rwl_21 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_22 wwl_22 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_22 rwl_22 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_23 wwl_23 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_23 rwl_23 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_24 wwl_24 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_24 rwl_24 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_25 wwl_25 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_25 rwl_25 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_26 wwl_26 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_26 rwl_26 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_27 wwl_27 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_27 rwl_27 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_28 wwl_28 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_28 rwl_28 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_29 wwl_29 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_29 rwl_29 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_30 wwl_30 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '0*vpp+1*vnn' 11.1e-9 '0*vpp+1*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_30 rwl_30 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '0*vdd+1*vss' 30.1e-9 '0*vdd+1*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vww_31 wwl_31 0 PWL(0 '0*vpp+1*vnn' 1e-9 '0*vpp+1*vnn' 1.1e-9 '1*vpp+0*vnn' 11.1e-9 '1*vpp+0*vnn' 11.2e-9 '0*vpp+1*vnn' 40e-9 '0*vpp+1*vnn')
vrw_31 rwl_31 0 PWL(0 '0*vdd+1*vss' 20e-9 '0*vdd+1*vss' 20.1e-9 '1*vdd+0*vss' 30.1e-9 '1*vdd+0*vss' 30.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vwb_0 wbl_0 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_0 rbl_0 0 DC='vss'
vwb_1 wbl_1 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_1 rbl_1 0 DC='vss'
vwb_2 wbl_2 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_2 rbl_2 0 DC='vss'
vwb_3 wbl_3 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_3 rbl_3 0 DC='vss'
vwb_4 wbl_4 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_4 rbl_4 0 DC='vss'
vwb_5 wbl_5 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_5 rbl_5 0 DC='vss'
vwb_6 wbl_6 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_6 rbl_6 0 DC='vss'
vwb_7 wbl_7 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_7 rbl_7 0 DC='vss'
vwb_8 wbl_8 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_8 rbl_8 0 DC='vss'
vwb_9 wbl_9 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_9 rbl_9 0 DC='vss'
vwb_10 wbl_10 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_10 rbl_10 0 DC='vss'
vwb_11 wbl_11 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_11 rbl_11 0 DC='vss'
vwb_12 wbl_12 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_12 rbl_12 0 DC='vss'
vwb_13 wbl_13 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_13 rbl_13 0 DC='vss'
vwb_14 wbl_14 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_14 rbl_14 0 DC='vss'
vwb_15 wbl_15 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_15 rbl_15 0 DC='vss'
vwb_16 wbl_16 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_16 rbl_16 0 DC='vss'
vwb_17 wbl_17 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_17 rbl_17 0 DC='vss'
vwb_18 wbl_18 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_18 rbl_18 0 DC='vss'
vwb_19 wbl_19 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_19 rbl_19 0 DC='vss'
vwb_20 wbl_20 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_20 rbl_20 0 DC='vss'
vwb_21 wbl_21 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_21 rbl_21 0 DC='vss'
vwb_22 wbl_22 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_22 rbl_22 0 DC='vss'
vwb_23 wbl_23 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_23 rbl_23 0 DC='vss'
vwb_24 wbl_24 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_24 rbl_24 0 DC='vss'
vwb_25 wbl_25 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_25 rbl_25 0 DC='vss'
vwb_26 wbl_26 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_26 rbl_26 0 DC='vss'
vwb_27 wbl_27 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_27 rbl_27 0 DC='vss'
vwb_28 wbl_28 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_28 rbl_28 0 DC='vss'
vwb_29 wbl_29 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_29 rbl_29 0 DC='vss'
vwb_30 wbl_30 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '0*vdd+1*vss' 12.1e-9 '0*vdd+1*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_30 rbl_30 0 DC='vss'
vwb_31 wbl_31 0 PWL(0 '0*vdd+1*vss' 1e-9 '0*vdd+1*vss' 1.1e-9 '1*vdd+0*vss' 12.1e-9 '1*vdd+0*vss' 12.2e-9 '0*vdd+1*vss' 40e-9 '0*vdd+1*vss')
vrb_31 rbl_31 0 DC='vss'
.TRAN 'timestep' 'sim_time'
vdd vdd 0 DC='vdd'
.END